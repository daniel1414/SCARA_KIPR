��   &��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����DMR_GRP_�T  � �$MA��R_DO�NE  $O�T_MINUS �  	GPL�N8COUNP �T REF>wPO�OtlTpBC�KLSH_SIG�oSEACHMS9T>pSPC�
��MOVB RADAPT_INERP ��FRIC�
C�OL_P M�
G�RAV��� HI9S��DSP?��HIFT_ERR-O�  �NAp�MCHY SwAR�M_PARA#� d7ANGC zM2pCLDE��CALIB� D~B$GEAR�=2� RING��< �PLCL*w ��STA� >mTRQ_M���LINK"2&SX�<*Y<*Z/)II*IzW*Ie$C�RV*� L $� E�NBpV_DEBuU��!PNU;%�� UNEVEox��!8� �$�A�SS  �����!����� V?IRTUAL�/1�' 1 5�� ��� ��b?M?�?q?�?@�?�?�?�?O�6��� A I�91HO6M��1 �� �����P��� G��5O�O1O [L�O�O�O�O�O_�KA_GR0_m__j_�_���d�_�_�_�_��=gL���_"o?�#o��@�Cohozo�o�o �o�o�o�o�o
.�_ 5YgwQ�4  2�_��� � ��$�6�H�Z���<���������̏ޏ�����&�8�J�����$% 15B1D�U5a���� �_���_�ϟ��,� �)�b�M���q����� ��ݯ�����(��L� 7�p�[�m�����ʿ�� �տ߯!��H�߿l� Wϐ�{ϴϟϱ����� ���2��#�e�'ߌ� #߰ߛ��߿������� .��R�=�v�]�gߩ� k���g�������<� '�9�r�]��������� ��������8#\ G�k}���� ����1�X�| g������� /	/B/)/3u/7/�/ 3/�/�/�/�/?�/?�>?)?b?M?�?[�RVk�r�`{?�?s?'  BVoKgx�?&O�8OJO\OnO�O�O�O � 6`
�  �:  R`�������������������������@$����\�����C���@�@����C��O_*_<_N_`_r_ �_�_�_�_�_�_�?o �_&o8oo\oO�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� Iof�Q���q�����so �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ����Տʯ���կ� ŏ"�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� �����������R� 9�v�)��߬߾����� ����*�<�N�`�r� ������������ �&�8�J�\�c߀�k� ������������" 4FXj|��� ����0B Tfx������ ��/�/>/��b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O+/HO3OlOSO�OC/ �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo}O�o�o