��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG  �D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!� ETH_�FLTR.� �$�   ��FTP_CTR�L. @� LOsG_8	CMO>�$DNLD_F�ILTE� � SUBDIRCAP"m� HO��NT.� 4� H�ZA?DDRTYP� A =H� NGTHph���z +LSP� D $ROB�OTIG cPEEyR�� MASKa�MRU~OMGD�EVl���RDM:*�DIS����TCPI�/ �3 $ARPSIyZoK_IPFp�W_MC-�F_�IN0FA~LAsSS�5HO_� �INFO��TEL� P�����R WORD � $ACCE�� LV�$TI�MEOUTuOR�T �ICEU�S�  � ��$O#  �����!��
��
� V?IRTUAL�/�!�'0 �%
�"��F��F��04+5��'�� =��!h�!j?����; x?�5�=y2~;#"SHAR� �19  Pf?O(4OHO7OlO /O�OSO�OwO�O�O�O _�O2_�OV__z_=_ �_a_s_�_�_�_�_o �_@ooovo9o�o]o �o�o�o�o�o< �o`#�G�k� ����&��J�� n�1�C���g�ȏ��� ���ӏ�F�	�j�-� ��Q���u����ן��ϟ0��7z _LIS�T 1�=x!�1.k�09��j�1|{��255.��Lr����05i�2p����砖�����̯ަ3 诂�_�� �2�D�ަ4`���װ��������ަ5ؿ��O����"�4�ަ6Pς���vψ��Ϭ� �$��Q>�$% =�/5+5�U�o!R��)��0H�!� ����r?j3_tpd��31� � �!!KC�� �߿�(�'6��!�C� ;�����!CON� ����=��smond���