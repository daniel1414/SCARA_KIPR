��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG�D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!  �ET�H_FLTR.�  $� �  �FTP�_CTRL. =@� LOG_8	�CMO>$DN�LD_FILTE�� � SUBDIR�CAP"� HOv��NT. 4� �H�ZADDRT�YP� A H� NG#THph��z +�LSP D $ROBOTIG �cPEER�� MwASKaMRU~�OMGDEVl�� RDM*�D�IS�� �OTCPI�/ 3 �$ARPSIZ�oK_IPFpW�_MC-�F_I�N0FA~LAS�S�5HO_� I�NFO��TEL�� P�����R WORD  $ACCE� �LV�$TIM�EOUTuORT� �ICEUS��    �$�O#  �����!��
��
� VIRTUAL�/�!'|0 �%
���F����04+5A�'�� =��!�!�j?����;� x?�5�=2�~;#"SHAR� 1}9  Pf?O(4OHO7OlO/O �OSO�OwO�O�O�O_ �O2_�OV__z_=_�_ a_s_�_�_�_�_o�_ @ooovo9o�o]o�o �o�o�o�o<�o `#�G�k�� ���&��J��n� 1�C���g�ȏ��쏯� �ӏ�F�	�j�-��� Q���u����ן�ϟ�0��7z _LIST� 1�=x!1E.k�09��j�1{�>�255.��r�&���05i�2p���@砖�����̯ަ3诀��_�� �2�D�ަ4 `���װ��������ަ5ؿ��O����"�4�ަ6Pς���vψϚό�� �$��Q>�$% =,8+5U��o!R��)��0H!�� ����rj�3_tpd��31 |� �!!KC� ��߿�(�'6��!�C� ;�����!�CON� �������smond���