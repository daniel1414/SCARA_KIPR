��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
� �A�PCOUPLED�1 $[PP_�PROCES0 �� �1�GP�CUREQ1 �� $SOFT�; T_ID�TO�TAL_EQ� �$,NO/PS�_SPI_IND�E��$DX�S�CREEN_NA�ME �SIGNj��&�PK_FI� �	$THKY�P�ANE7  	�$DUMMY12*� �3�4�G�RG_STR1� � $TIT^�$I��1&@�$�$�$5&U6&7&8&9'0''�%!'�%�5'1?'1I'1S'1�]'2h"GSBN_�CFG1  8� $CNV_J�NT_* �DAT�A_CMNT�!?$FLAGSL*�CHECK��A�T_CELLSE�TUP  P�� HOME_IO�� %:3MAC{ROF2REPRO8^�DRUNCD��i2SMp5H UTO�BACKU0 �� �	DEVI�C#TIh�$5DFD�ST�0�B 3$INTER�VAL�DISP�_UNIT��0_�DO�6ERR�9FgR_Fa�IN�GRES�!Y0Qy_�3t4C_WA�4H�12HGW~0�$	Y �$DB� � CO5MqW�MOJWH�.
 \�VE��1$F �A��$O��D�B�CTM�P1_F�E2�G1Q_�3�B�2GX_�D�# d �$CARD_EX�IST�$FS?SB_TYPitA?HKBD_S�B�1�AGN G� �$SLOT_NUyMZIQPREV���G �1_EDI}T1 � h1�G=H0S?@f%�$EPY$O�Pc �0LEToE_OKRUS�oP_CRQ$�4x�VAZ0LACIw�Y1�R@Pk �1w@M{ENP$D�V��Q�P��A��nQLv*OUyR ,lA��0V1AB0~ O�L]eR"2CAM_�;1 x�f$ATTR�MP0�ANN�@�IMG?_HEIGHQ�c�WIDTH�VT�C�U�0F_ASwPECQ$M@gEXP;�@AX�f��CFT X O$GR� � S!1z�@B`NFLI�`<t
UIREs3��tGITCH~C�`N�.0S�d_L�`�CL�"�`EDkp;tL0J*DS�0>0�zra�!�hp;G0 � 
$WARNM'@�f�+P� �s�pNS=T� CORN��1�FLTR�uTRA�T@0T�p  $ACC�1
� ���ORI	`!S<{�RTq0_S�B�qHuGI1 [ �Tpu3I8�TYPVD+P*2 �`v@�� 1R*HD�cJ�* ���2��3��4���5��6��7��8���9�mQCO�$ <� #5x�s1�v`O_M�@�C �t 0Ev�NG��ABA� �c��@YQ������@������P�0����x�p�PyP�2� h����J�_R���BC�J��2�J	VP�CR��}@w��lu�tP_}0OF� �2  @� RO_�����aIT8C��N'OM_�0�1åq384 ��T �#�d��@xP��J}EX��G�0� .��p�
�$TF`��C$MDM3��TO�3&@U=0^�� �H�2J�C1{�E͡� vE��uF�uF��0CPho@�a� 	P$@`�PU�3�f)�"��)�AX 1rDU�6�$AI�3BUFpV��o@�! |�plڶ�pPI��PZ�MY�Mf�̰i�}FZ�SIMQS���/��A-����jx Tp{zM��P�B^�FACTqbGPEW6��Ҡ��v��[MCc� �$}1�JB�p;�}1DEC�Gڙ�G��A-�b� �ě0CHNS_E;MP��$GO���B+P_��q3�p�@Pۤ��TC��{r��q0�s ��a�/�� �B���!	����JR!0��SEGKFR��Iv �aR��TjpN%S+�PVF�����ʹY�K����a1�)B���( 'j�Av�u�ct� �aD�.0���*�LQ��D�SIZC�������T��O�����aRSINF�����jq�� C��C����LW������x�CRCLuFCCCkpy�����N}�� �bA�������d��DwIC��C���r��`+ P��z�2EV2��zFH_��FpN�t/�>�����H�1Q��!  � ��Qx����U�kp�2@ ��a��s�+���q}RT!x "� 4�4u2��tAR���`�CW�$LG�p��B@�1�Pr�P�t�aA?@�z�ϣ~0R�ӲM�E�`8�oC�RAs3�AZ����pb��OS�FC�b�`�`F�Mp�� �0��ADI S+�aV%��b�z��p E$�pRp�cV�S�P�L�a+QMP5�`Y8C���Me�pU��aU�S" $=�TIT�1�S�SG1��#�8��DBPXWO! zT#��$SK���FDBTmTRLS$l�Q0TQ��P`�P�D�q�1LAY_CAL�1�R^0o f7#PL)A�Q�D'a�73a�7��)2!S�%2?�PRj� �
*0���S& l=�A$��$ �
*�L�9'�?'�U�T)(ODCS)#ODgENE��*BO�'Ӳ0RE�pB+�H �Ou�&$L�C'$�3R�h�K2�LVO�_D~!U�ROSbrq�v�R�����CRIGGER��FPA�S��6�ET�URN�B�cMR_�}�TUbp���@EkWM$���GN=`����BLA��TUܡ�($P�)$PD s�*hP3a��C�TΣ@DO>���D�A����FGO_AWA�Y�BMO"�a�!�*0CS_P,<aISt�� �� �s �S#�Q���Rw� cV��Qw2�VW��'d'NTV(��RV;��@��~��mgŃ��Jtx��<@��SAFEڥ�f_SV�bEXC�LUT��� ON�L���cYfЀ�y�O{TEuHI_V} >��PPLY_�q7��VRFY_b3 ��Sj L�_ -�h@0��_y�1� �(2�PSG�  .�rŐ1PNQ5�� _q���;P��Vby|rsvANNUN<@�$�tKIDX�UR�c[P�� �y�qi �z�v�2E�F�PI<B/��$1F�r�$АOTQP�A� $DUMMAY��&���&���*0|t�U0 `  �HE�\���^r�cYR�r SUFFI��A�Pa0��P)�5#�u6#�N)1MSW�U�1 8��KEYI��4�TM�A��ځ3QFՆINݱv�JDj �P2 D��HOST�0!������`�������EM&�����*0SBL� UL��3 Z����D�*0T�@S4 �� $���USAMPa༥.������V �I�@��$SUB����;@c����3��SAV�������`����`�vP$�@yEC!	0YN_B375 0��DI�t�P�O\�M��#$E�R�_IB� �ENOC2_S�T6X��2������ �cG���0 S72��1��A�����8   ��Ǜ��@PK�Dk!<uq��AVERҁ������DSP�ܢPC?���26�\�����oVALU�HE ��M_�IP(�ܣOkPP� 5�THЈ�ͫ��S` 4�.�F�B�6d��~�� 5�SiC?q���ET��9ȂFULL_DU���qKP�ԝ������OT�"�QPN_OAUTOS:�C$YĪ�Z� ���*X�C��h�CE26���V�L� ;/H *h�L� �����$P��wc�� �1�Ʃ1��C��Ƨ���T����7��8��9�ʩ0����1��1��1�	�1�1#�10�1*=�1J�2X�2����U2��2	�2�2#�U20�2=�2J�3Xڥ3��3����3	�3��3#�30�3=�3�J�4X����SE�2< <8�Z�����I��e�$�}Ń�FqE5P?PT= ,f���a? �P�?Qi��e�i�E�P�q�(1aT>F��$TP$!$VA�RI����UP2f1p? 7���TD��@s��p��������wBAC2@ T� ���$uP�*��Þ0� IFIw�0�P� � *)PB"��F0P�>TAt ;u�"�"pu STvt: @�bt�@�l�6	sC2	>0���S����/bF��FOR�CEUPsr��FL+US�pHfNn����bD_CM�PE8v*IN_t�\e`�REM� F�a��a�0�Te�KrdN~�eEFF��j�PINJa�OV�M�OVA�TR3OV��DT	��DTMX,A��P *��0M(xR#�0�CL*_��u*�Pr�2{_XЉ_T�+*X��PASaD% ��(װ�1`�&_A@�RQ�LIMIT�_�4�� M��C9L�tˑRIVW�n*2EAR�IOx#PC�P���B�R�cCMQP*�b !�GCLF�#�1DY��8} �q�35T�%D�G���0�5�#pFsSSt0��B P�(�1�A��`_�1�8J�11��E�C�13 K=5 F�GRA��g�C��k�`W�OyN��"EBUGwc�tBxJpC ��_E �D ��K� _�TERM�EE�EN�AORIS�@F�E
�SM_�`����@G�EP��TAr�IH�EcP�UP���I� -�Q���D|`�C|PE$SE�G#Z�0EL�eUS]E�PNFIzLR�T�kA,��DTF$U9F�`O�$\��aD�P/���Wi@T���t �cNSTTPA�T��h��RPTHJKa-�E
�65MR<p&� WUw�&�Q�LQR<`�Y�qSHFT��MQ�Q>�X_SHOR�*�J�F �@$�GM`H��u OVRq��q6`I�`4U� �aAY#LO���"J�Iu2b�p�Q��oƸ�ERV�� �a� 6j�WnP�R~�PE �e��E Rb1PpŏASYM|�p�MQWJ`W�� E���Qy�b0�U7tnPI��Uw��/�ePo��`o�fgO�RnPM�G@SkMTfJg�GR��aC�qPA|P��p=���K � FNTOCFQ�P9`N $OP@/��(#��N �!O�ڐKRE
�RdS�QO��,��Re�R�UN��%�a#e$PWRf0IM@��bR_ ����=�mR LVBH|�_ADDR$�?H_LENG�Rǁ����T�R� SO�M H�S���~��`������	�SE!�u���S:�MN�1N��p��F���OL��8�3�3�=��ACROc�z�P�$��[·a;�  �OSUP���r_�I���q�q1�ѭʓ��ԙ X!՘Y1՘t!՘	�ԙ�лE"IO���D�ϗA�ߕ9�gO �$���p)_OFF�b�;�PRM_Ò��qTTP_[�H�jP (��OBJ؍2��#$$�LE�S���Q � ����AB_�!Tġ��S�p;x LV朳KR32@�HIT�COUBGE�LOہ磴!��@���"�G#�SS��HQWD�SQjR�lp�INCPU4BVISIO�����Ğ�
�����	� �IO�LNS� 0C^$SL�r@oPUT_�$@���PV0�ɱ)F_�AS�2T $L   �� =a0U�@9`�dQٵ��䳊`HY�#�]�6����UO�3U `"�{�$�@5"M�5 Tƥ�R�P;�@��ǿ�T��µƑ�UeJeV]���NEfg�JOG{W��DIS���K��� �3W �XХQVv��P;�CTyR�S:�FLAGBBv�LG�tX �� ����aCLG_SIZ����d �����FD��I�اؓ�� �ث@�֎����	�d  	��	��	�@	�% SCH_��R���aBRg�Nє�Y��!AE�2��p�J U}��}��pL��|�DAU��EA�����t����GH�rt�%�BOO>Zh A<�f0�IT2���@8�REC�SCRB�=��D:�����MARG �<18��0��a�%�Sȣ$�W?�%����0�JGM��MNC�Hz%�FNKEY���K��PRG��UqF��g`��FWD���HL	STP��V`��mP������RS;	Hp��-�Cid6r0�.0s��	U|���r� Xb��P�E���G��`CPO�
.�M��FOCU�RGE]X,�TUI��I��p�K|�V��V�� ��A`B���p�A`�9Nu��SANA%�FRޚ�VAILy�CL�P1uDCS_HIyD�
��O�X1��S� ��S�V�I�GN��~�ӽ�\�Tx��0%�BUFF�1�[5�o`T�$ ��� ����B����A��\5�o`ܰ��\c��pOS1�%2�%�3�!�$��0] � ܩ�qEU���.��IDX�tP�bD�aO� ��Q6ST|��R��YV�@1 \$EO6CO;�{��^6q6L�%��0^ L��K�[@`�9`(���S���:�����x��_ _ o�p�ÐЌ�� C�@Cp�` =�� CLDP|�uTRQLI��Ft
�4I"DFLGV�"@1�VC�D)�VGr�LD8VE@DVEORG
�q iB_�g�H
��d�D�ta �M�@Dr1D
VES�pT4@I��@T}VRCLMC%T`�O�O7Y���MI�έtb dy��!RQzI�M�DSTB��0 �VO�XAX�r �X�\EXC#ES6��!vRM_��q%c�0�RtsU<�j�pd��V_A�Z���(k�_�X@K�te� \����/�$MB�s�LI���cREQUIR�b��l���hODEBU��sQL�0M,�f�r=��`�����%R	bND���p�pg0w�n�?�sDC��IN����p�,x' �NV���K��eP�ST� h��L�OC�&RI���%E�X�vÀ�!�QsQOwDAQ,�i X��3ON���MF\��� �v9�2%��5�uk�0�� �FX�PIGG>�� j �M��2�!���3��4R �%?3;�|�K�|�Z�G`�E�DATA{'��E��U��b"���NZ"k t $MD��I��)Ɔ ф��ф�H�p�`Ѕ�X�҃ANSWe�ф�!'х�D[�)�r��P��l[ �PCU��V��X@�uRR2��m �D���a���Rd$C'ALI�P"�G�w��2��RIN��z�<Nu�NTEڰ�"nI�`��°r��ڰ_N���oÕޒi�oT۔bpn�DIVmVDH�Ptݐ��q� $V���+s1$��$Z �"��� �"f�_�e��rH �$BE�LT>��1ACCE�L!������IR!C��P��t�T31h�$PS�P'B�0���Ȧ<C���������P�ATH������3ТZ��Q_�!U�2�8��R� C堌�_MGP�$DDU���/�$FWh�����q�ء���f�DE��PP�ABNاROTS�PEEH��!��4@J���!��P���$OUSE_���P��FO�SY��g�Q B��YNyPAO��OF�F��MOUR�N�G�O�OL�L�INC.��q��u��Rn�<PP�RENCS����`�Rȡ���TŠIN'2�IТ���`R�VE�S�{���23_UP�I���LOWL! � �4@���D� �R {`���0��5bCΐ��gMOS4 LdMO����PWPERCH   �OV��b��! m�@1�^T@1�s��hP�`�� V5�'`ѡ���L���Ig����U�P�Ӛ���TRK|v�#2AYLOAA ��$a1�Т@�5�p40���RTI(a|�40MO����R$b�@N��T���w�L���"f�D�UM2,�S_BC?KLSH_CТ�� B�A�u�'�Y������x6�x�aQCLALz ����Ar�`�CHKt4@+5SH�RTY S��}%�A��_:36�'_UM(`n�C{�c��SCL��ʰLMT�_J1_LS��P������E�������8������SPC��;����	��PCsѦ�H��0�`Y�q�C3P�2X�Tc�g�CN_��N���i��SH ���V 	�*3�Ň�=Т�AC� y�SH:3��g� �ƝA���s�4�ѡ̬�c�PAx�l�_Pw�[�_5@��8�V�4AH�ZK�JGG"M���OG[��TORQU��ON.�Q靰wb0LҠᝰ�_W��1�_A��G��M��I*�I�IM�F�p�aJPQ2(�A_�VC��0�T�RS"1Y.�Pm/�R`%JRKY,�"�&~PDBL_SMh�:RM)p_DLG�RGRV��$G��$M���!H_ �#�:CcOS;`�8LN�  ;;\%B4G�=9M�=9!y:g<-!�%Z60L־!cMYD1�8$2TH*=��9THET0�N�K23M�BA�E0C-BFCBA�C�Q�R�,B$:AG�:AFSB8G�XBEGTSaʱC��qW4&�Dg3<�Gv3$DUH�Ih��Aw�x��R�F���QQ����v$NEd�I F0Y�`R�E��$%��1�A�5#U,W
581LCPH(eR��RS\% tSg5tSv5R�6�S�Z�6%�VEXV:X7�]\UVlZVy[V�[V�[UV�[V�[V�YHEX@^Vdb\]�{hy[H�[UH�[H�[H�[H�Y�O6\OEXO�i[^O�lZOy[O�[O�[O*�[O�[O�6FR'A��yg5�t8WSPBA?LANCE_�1�s�LEo@H_�5SP���X6�rg6�rv6PFULC�x��w�v5�Ț1n}�UTO_<C�nT1T2G���2N*�z���g���k���@ע����T��O�����INSEGz�%�REV��%���gDIF��1o҇6�1p�@OBȁ��#��MI��5��$L�CHWAR����A�B*y�$MEC�H0A�0>�D�Y�AX�>�P��]�W(�<�q� 
^������RO�BV�CR�Ҡ�RJ���MSK_�pj�s� P R�_��R ��H�Ҕ��1����ԲҐ����Ґ&�IN����MTCOM�_CD n�t  �P�ڀ��$NO�RE��9���(�7u 8�GR�I��SD�@ABJ�$?XYZ_DA9Q���DEBU��M���U�v �p$�COD�� ��o�J��j�$BUFI�NDX԰����M{ORœw $1��U��-��v�F����ѣ�Gܢx � $SIMULXૠ���$���OBJ�E�p$�ADJUS<B�5�AY_Io���Dc����G�_FIJ�=�T����� ����������Հ�P:��D�FRI��׵MT��RO���E�<���OPWO� ɐ�y0��SYSByU�PΠ$SOP�ȼ�#�'�U&�ՀPR�UN�M�PA�DpL�H�!���_OU�!�A���r�$��I�MAG��ϐ�@Pf��IM����IN� �u£�RGOVRD̱>°Ѐ�P����԰�@L_:����m� SRB� �@M���EDՠJ� ��N�pM.������SL��pɐz x $�OVSL��SDI��DEXqk�i�=!H{��Ѕ�V���N�р�{��Њӟךط�M��!t G�_SsET�ɐ{ @����g���RI&���
B��_4A��	������ׁ@��  | HxϑI�J�ATUS��$TRC�@ǰˢND�BTMM�7�Ij����4��#�,�ɐ} DϐE~�k�A�`�EۂBᏱ
��B�EXEH�Z�ќ��{�b��~��АG�UP���$����XNN�m�=!p�L!p� �P�G&��!UB�6�g��6�
�JMP�WAI� P��N�L�O��1�F��#�$�RCVFAIL_C�1�Q�R��Q�Z��M� 𣕠���0R_{PL
�DBTBm��1�BWD��A�UM���IGe���m��� TNL� ����R���.�Ep�һ��!�DEFSPy� �� Lϐd�7 _8: H�HUNI��r��F ��R��^�� _L*��P@��P�ȑ����F����Ѐ��p:��N�pKET�}��� P��ȑ� h~W�ARSIZE���l���S@�OR~
�FORMAT3����COJ����EM2V�lUX���� �PLI��ȑ� � $#�P_S�WI�i���AX�����AL_ ���E A��B�,@C���Dj�$E����uC_��	� � � ���q�J3�@����TIA�4�5�6��MOM�������#�Be�AD�&�&6�PU;@NR�J%��J%�7EŔ�?� A$PI�F� ޑ��$�%�#�%�#�% =D�&�+QD�DpсF����U���g�SPEED�`Gd*4f�7 167f���16g3@8p��O9��f�SAM�p�맣417�3f�MOV ���D�1ƀ�E�4�E�17 1��42��������5n��Hm��3IN2Ln�39HUK0Df��;J{HRD{K�KGAM�M�v�A�$GE�T��ȠL�D� �
�b�LIBR��I.��$HI��_��P�$�bVE�XA^:P+VLW]XVO\:Y|V�+V�V����� $PDCK�DU�L�_�0�� �.B �m!E�W��T&�Y~r �$I�RS�D��&����(�LE�ޑ�Oh�)`���H�ɐ�P~��UR_SCR����a^��S_SAV�E_D�īe��NO�C����`�D� �&�i��)�iapz{ p���&Ex@�q��0 �B���5G�2�+8!� ;6��g8�w�ucs�1��tiHM{%� �� ��!G����c�w���`�ζ�qW�`��$�� 0�N ��R�qM��H��CLG�GM�aǒ� � $PYr��$Ww�+�NG t��w��u��u�� u��������@[L�JnX� O�mZ��8GQ�Ŕ� pW�#�c�&�o�o#5t��_)�� |W� ��`��������`�ޗɖ�EQ��Eϡ(F���b�Ϡ����P��PM��QU��0 � 8� Q�COUa1�QTHHOL��QHY�SES�1[�UE�G��b� OM�  b�P4�U�UNI�.J� �O��)�� P�������a��ROG�j��2���O𤥥c�󠉠IwNFO(�� ��hث�
��1OI��� (`SLEQ�"6D�5D�ܦ����D$S𿠒��VPO�P�0j#3QEMPNU��Ύ�AUT�a��CO�PY�1�಼��`M"��N������CT��} �RGADJ(�e��X#�_$� ('��'�W%�P%�]`�'�:3�;�EX��Y%C��1@OՐ(����_NA�1�!S���i����M�� � ��p�P�OR��Ì&��SReV��)����DIT_p��� ��
��
�w�
�5�6�7��8��1S�b������MC_Fe�B�pL�a�a�;�Rq� ���/��җ#�0��k�n�� ,`FL��L��`YN{���Mp�=C��PWR���z�����DELA ���6Y�ADR��� ��QSKIP{%�� �����OŀNT2�1�0*�P_���� I�`߂̐`��#`�3 `��n�kn�;�m�HРm�U�m�b�m�98a��J2R.0��� 46� EX�@TQ�� ��q����������y`RDCx�� ���X��RF�E@A�Y�_�X�DRGEA�R_�@IO�t=bF�LG���EPC���UM_���J�2TH2N�# � �1�UA�G�@TN�P �"���M���-�I���4�REF:�11(�� l!��ENAB� ��TPE2`{� 8Wܠ� M�q�CL��R�w��2'�-?QPcu��3'��@�����4'�'9K]o��5'��������6'�!/3/E/�W/i/{/ @�!7'��/�/�/�/�/�/
�8'�?-???Q?xc?u?�SMSK(������ E�a~�qREMOTE���
��`/B`��q&-CIO�UQEI�0��R� W\`��� �/���-�����ҿ����ՈB$DSB_S�IGN'a�q����C���pS232�3E���$�DEVI�CEUSKC�r�rP�ARIT!�AOP�BIT�q��OWCONTR���q��0�rCUPM�sU_XTASK�SNq���P�DTATU�p��C3`���u�e�_��pC��$FRE?EFROMS����Θ�GETA`��UPeD��AEbSPTP����� !�8$USA�����9h�{�ERIO���`Ր�RY�U�B_�`��P8�QQfWRK�?�<�Dh�3fh��6FRI�END�qg�$U�F�U�p`TOOL�wfMYd�$LENGTH_VTߤ�FIR��cM�SE<�@�iUFINtrа�ARGIaF�A'ITIi�gXF�i6�fG2�WG1�� �Sr$wPR��sau��O_�@�P��xQRE`���SU�ءTC�8N�=qyv�G��]R
���u��Q�A��hz hZUz�ZU�t���{P>�T�X �P��L��TcH��hh�(U�T�SG��WX�)�	�r>�D���.��`C�z�N�b��$�v 2�!�-a' 3i�1?h.`21k2��31k3?j���@i���`�6{��s{��r$V�J�bV�eV���a �qYr���O�[V{�@���hv3Ru�^pib��P5S��E�$���c��5$A8й�P!R)��u,�S���@p���D�Q�¯ 0pD�v���P�N����!�P�P>p ��
�USzA/� �\�R��GA�_�Š��Ny@AXQ��Ag`L�ag�p�/THIC'a��-����QTFE���m��IF_CH'cp�I0_����6D�G1՘٤�*��h��`��_J�F�PRW�I��R�VATF�� �`\�'�f`��)�DO�e�)�COUW�C�AX�I�D�OFFSEZ�TRIG�sz�,�@)�#g���z�H��<��g�IGMA�P�a�\���ȸORG_�UNEV#@Ͳ ��SD���d ��$����GROU[A�TOa�Q�wDSP#�JOGV�LS8�_PV�3RO��p�U�mpEVKEP��#IR?�_�=pM ���AP���E��������SYSv��B��PG��BRKYr����b�\��������k��ADVQ�y�BSO�C�C@N�DUM�MY14��`SV��DE_OP1SS�FSPD_OVR����C~�N�Q�OIR\׶0N�P]�F��l]�<�OV?�SF��a����F���Ac�As��؁a�BLCHDL>�RECOVM��P�<�W�`M<��?�R�O1S�K�_a�_�s @���`VERt��$OFS�`CV�@_bWDv� �r��X�R��9�TR%QA��E_FDO��MOB_CM[A��B/��BLl�_¦�l��V@�qDb�P����G����AM�Ú�yP��'��_M��>R��HC4�8$CA2���Ȱ��8$HBK�Q��N�IO1e]�iAA�PPAQ�}�b���u���iB4�DVC_DB �c�񓡦B����A���1��'���3��-�ATIO�@��FPM�qUDc1�HFCABH� 0bFs�p�p��Ea<��_BP��SUBCP	Uk�I�S%��@���䀬P�s�,���B��$HW_C!��i���x�A'q\�l$U�NIT��l�AT�}����I�CYCL���NECA#��F�LTR_2_FI`Ҥ�H)�FEaLPU˼����_SCTosF�_�F��
v�
FqS�A���CHAJa�^���3R�RSD�1�B ё�l�i@_T���PRO ~�)PE%M�0_���8�3�� �<�*%DI��P��RAILAC4��rM��LOГc+�i���-��-'�+PR��S{q*��!�C���@	&�FUN9C�³�RIN�pZ�0+`? �$(QRA� mr� 9��#��G��#W3AR�:�BLuq�'�4A;88DA`���!I835LD�P A�A�q3h��!��q3�TI���5�β�pR�IA�Q�BAF� P �A���1��5��T����EMJ�I1Q��DFa_�`�ӨQ��LMt�{FA�`HRDYd�P�`RSoq+`Q0>EMULSE�`��<�E� ���I������$]a$6�Q$�Q�,���� x��EaG�P�AРAAR�2)�09mb�E50��wAXE&�ROB#��W�ac�_�M�SY����Ae�VSWWR�ذ�M12�� STR�"Ņ�d�h�E� !	CUq#��lqBhP3�oV��)��OT�Pv� 	$�ARYg�ЦR_!�`	T�FI���j�$LINK(�1w��Q�_eS3��CU��RXYZ@Q��[��	co��Q�RJ�X�PB!��"Kd0�
 � LcFIeg`3�D�9Ԫ$<�_JN�p"�e��SA�OP_~T2�[53�NqTB�aNB2�bC9��DUQ�BV=6r%TURNb����u�Q�!h�?�gFL�)���B�@+pekZ7�3�I� 1�nPKH�M��BV8r%����c�ORQ&�!�# mX�C�����갦��up��.�<��tOVE�q��Mj�tC�zC��B�W�Fq�� � ��� j�0���qw�P� ���	��q���zC��L5��!ERM��!	v"!E8P���#؄A���id�%"�WP1MP1AX�bP1��&!�Q2� 2!>�\A>���=��`=� p=�ep=��p=��@=� JQ=�@:�@J�@Z� @j�@z�@��@���@��@��ב˙DEBU�$�!�1($�{�P��R�g� � AB�P'N�[��sVְ� 
����Ϥ��Ϥ aڧ$aڧ�aڧqڧ eqڧ�qڧ�A�4�`�2\�RLcLABbb�u�� ���1sE� �E�R�9P � $�8`� A�!��P�OB�FЉ�P����_�MRA��� d �O0T<�\�ERR�:�2�0TY�aI�A�Vb`,���TOQ�+�i�L�@,�7R�􌴇 C�A � �p�T�P��< _VA1ْ.�V�2#c�2\�!2k�ȱ��op�ˠȱ�u�$W��6�V�A���$�"�0�,���6�Q�	��HE�LL_CFG�A�� 5e B_BAS��SR��p�� �CS��1�U1��%�22�32�U42�52�62�72�82��RO �8��Pf,`NLzA�cAB��H �ACK��>�i����`�`G@���_P�Ur�CO�@��OU��P0�W!��3�7�LTPX�_KAR����RE��&@P8 W1�0QUE� ��p9CCSTOPI_AL�����PU#p�Д���PSEM�d��M���TY��3SO��W�DI��p��}�L�1_TM��MANRQ��PE�ZV�$KEYSWITCHU#8���CHE9BEAT4!�!E�@LE�$
f�U4�F��5�K��_O_HOM�0O�#7REF�pPR�!)(�AUP��C��Op�0�ECOư_1`_I�OCM�d���m� �@��g�@� DH�Q� U۲{�Mw2xQ��p�cFORC�f3 4���OM�@ � @���3�U[SP�@1��$�@�3�4�1��NP�X_AS�¼ 0��ADD' h�$�SIZ�$VA�R2�D@TIP���� Ah�аJ�萲 �� �BS��AC<��%FRIFa��aSe�w	��NF򸍰Џ@� x�S�I�TEFsj"esSKGL}T�R7p&A����#P~STMTdJ�P�@;VBW�p�SHOW�R���SV
@�D�� �ԱA005pЁ " � '� '� '� 'U5)6)7)8)9)A)�@'v 'V�	&r`'F(JP�( )�P�(,)#`�(F)p��(`)�p�(z)1�)1��)1�)1�)1�)1��)2)2)2)2�,)29)2F)2S)2�`)2m)2z)2�)2��)2�)2�)2�)2��)3)3)3)3�,)39)3F)3S)3�`)3m)3z)3�)3��)3�)3�)3�)3��)4uI4)4)4�,)49)4F)4S)4�`)4m)4z)4�)4��)4�)4�)4�)4��)5uI5)5)5�,)59)5F)5S)5�`)5m)5z)5�)5��)5�)5�)5�)5��)6uI6)6)6�,)69)6F)6S)6�`)6m)6z)6�)6��)6�)6�)6�)6��)7uI7)7)7�,)79)7F)7S)7�`)7m)7z)7�)7��)7�)7�)7�)7��$��VPd�UP}D��  ����)�
 YSLO>��� � ��0�Q��TA�����ALU������CUT��F��ID�_L��HI�I~V$FILE_�?�+�$�󍰢�S�A��� hҰk�E_BLCKh�x��>��D_CPU���  ��� �B�T�b�q�	��R �G�
PWll�� �LA1�S������RUN u������8�u�?����?�� �T?�A�CC��X ;-$f�LEN��s����f�����I�J�L�OW_AXIh�F)1f�,�2��M��	�G�_��I��Y�8�թGTORn�f��D��<ܣ\LACE��Y�pf�ٳY��_MA� p��3�	�3�TCV:�[�	�T�\�{�q�| ������	���J���ŉMĴ�J9�����	�r�2�Ц��������ΠJK�VKо�#���#�3�J0l8�'�JJ/�JJ7�AAL'�]�/�]�W�e4X�5��{�N1��P��M�I�ڤLӠ_����b���� `u�GROU����}Bd NFLIC���REQUIRE��EBU��b�Ŷ��2�c�	�a�� ��� \APKPR�C �ܠ
a�;EN\�CLO��lهS_M`������
�a��� �F M�C6�{�����_MGV��C�l��؎�5����BRK��NOL������R�_LI��������J��P _��/��7��{��D���6L�O�8����>��� �ҍ�z��燡��PATH�������ᒨh��� $��ͰCN���CA �]���INFe�UC٠��%�C��UM.�Y��4���Ez�P���P�7�P�AYLOA�J2=L��R_ANE���L���������R_F2LSHRC��LO��$���2���>2�ACRL_�"�� �����H�b��$H��CFLEX�_�a�Je�� :r���	�t������	�������F1 ���ïկ�����E'�9�K�]�o� ���������$��г �#(ؿ�����	TR'�X ˲�` H��%�&�8�J�\� `�i�W�{ńϖϨϺ����J��� � `������ʁ��ATl�ðELt �5j�J����JE��gCTR�TN"�F�6	�HAND_�VB�_����� $f F2�֋���SWy3`������ $$M���R �ӅH�ѕL��E:�F�A�������I��A(��݀��A��A	��@��۪���D��D	�P2��G	�qYST��yQ4��yQN�DY �Z� �ּD�E��)�����������H$� � �P T�]�f�o�x����}3>�� {@`���n�vf��o�ASYM$������Ͱ����_SH��#�=� '��dLHG�Y�k�}���J��G��gs]y��_VI/C�x�ӵpV_UNI���t�#��J��re�r���t ���t�ð	G�(H:j��#PX��2A�H��N��EB��3EN/@��DI	�W#�O��e ^ ����S� � �BI�aAK� ���吂��U��0`�|�n�� � ]AME\?0�g��aT��PTpi0��5�����K�,p:�U�I��TKp�� $D�UMMY1�!$7PS_RF� i@k$��͑LA���YPV#��=�$GLB_T~@��ŕ5�ఁ`�CAӁ� XXI�	נ�STȱ��SBR��M21_�Vɲ8$SV_E�R��O��#�CLߐ�AuO炔��0�O� � D �ĐOB���3LO �f�S�y�ÐS�p�1wSYSS�ADR�1ܔ�5�TCH�@ �� ,f L���W_NA
����y5�SR>��l }J�J���F��B ���G���I���ID��� D���D���V�p�KYV� ��bu���ݻ�������);MtɁXSCSREi�W��E@�3ST��F�}��a¦Ǥ��0_�0AV�� TI�&����1�%������1���Z��O�PIS�1������UEЄ� ��񪠞�SG��1RS�M_����UNEX�CEP��ј�S_ ߑ��7��&�9�T���COU\ғ� �1֤�UE���؂6�y�PROGM�@FL�1$CU�&�PO�>��I_��H�� � 8\E��_HE_�������RY ?��0���������OU}S � @��~D�$BUTT/��R����COLUMx0��s�SERV�3���PANE�0V��:�TpGEUA|��F��ʡ)$HELyP��bETER5�)��E���Oq��30�� ;0��M`��U`��]`��SIN��-�TpNp���0�131� ��i�LN��ܓ �0���_����s$H_�0TEX�3�j�^�~$RELVB"D��~Ӑ�b���Ms�?,��p��4������#��USRVwIEWV�� <����U"�]@NFI<�0��FOCUA���7PRIx0m��h�� TRIP��m��UN��Є� x�`/��WARN�����SRTOL���&�Rs�O�cOR�NsRAUW�vT��	���VI�υ�� $��PA�TH���CACH�V#LOG��LI�M�r�S��BR'HwOSTǢ!�z��R|�OBOTƣV#IM� ��Si@��0r�������V�CPU_AVAIYL���EX�!�aN��} ~�Ma�Ua��]a ����{0�$BACKLAS�� �!�$"W��  �CT%s�@$T�OOLǤ$�_J;MP�� ����$SS�v4��V�SHIF`у�APB���ǤЇ�Rk(^�OSUR�3WRADI�$��_ ���%�м1�ぺ��$�LU�q$OUT?PUT_BM��IM���b� }p���#wTIL�'SCO�"�#C���$N�&N�' N6N7N#8���!u%=,�2�P#��`Є�<��DJU�rU��P�WAIT����<��:%0N�E~��YBOW� �� $��춤��SB"ITPEo�NEC/,B@D(D�PJǐp�Rv hE(��#=@�0�B�E/�M �KT���"y�� An�v!�OP�
MAS��W_DOآ�qT���D]����C��RD�ELAY��SJO �"X֡�c'T�3��``� ��,l�y�Y_�Ry�wR�#ƢA�?� 
��ZABC�� ��Rz��
���$$C�>X����Q��x���P�PVIRT��_�PABS�!��1� �U� < �Q (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П������*�<�K�`�AXgLMTZK��c7  �]�INf�x��\�PRE�Nk������LARMRE?COV �Y������@F �U/�QdK�� "�4�F�T���w�����<����, 
#o忶W�NGu k	? A   �,˾`PPLICu�?��U����Handling�Tool m� �
V7.70P/�36+��
��_3SWr�F0���� 43�ˊ�yϋ7DA7�철�
f��rm�N�one����O�հ�P�T���<�_+�V��R�v�7�UTO�RX l����n�HGAPON��Pe� an�U' D ;1�� �и������T�n�� Q 1M�  ��������	7�H嵡]��R��R ��a�,�H��B�?HTTHKYV��R �+�=�O������3� ���!�?�E�W�i�{� ����������/�� ;ASew�� ���+�7 =Oas���� �'/�//3/9/K/ ]/o/�/�/�/�/�/#? �/�/?/?5?G?Y?k? }?�?�?�?�?O�?�? O+O1OCOUOgOyO�O �O�O�O_�O�O	_'_ -_?_Q_c_u_�_�_�_ �_o�_�_o#o)o;o Mo_oqo�o�o�o�o �o�o%7I[ m������`��!�[���TO��C�U�DO_CLE�AN��5Ի�NM  	�Կ��+��=�O���_DSPDgRYR��HIa��@����ϟ��� �)�;�M�_�q�������MAX@���[����׳�X�����҂�7�PLUGG�У��ӮS�PRCt�B�"�������O�}�^5�SEGF{�KY� k�v������Ͽ��8�=�p�LAP���� o�Y�k�}Ϗϡϳ��π��������1�v�T�OTALզ��v�U�SENU���� ����ߎ���RG_S�TRING 1~s�
�Ml��S3�
��_ITwEM1��  n3� �����"�4�F�X�j� |���������������0�B�I/�O SIGNAL���Tryou�t Mode���Inp��Simu�lated��O�ut��OVE�RR�� = 10�0��In cy�cl����Pro?g Abor�����~�Status���	Heartb�eat��MH �FaulAler%	U�CUgy������� ���۞����6H Zl~����� ��/ /2/D/V/h/z/�WORy��۲! &�/�/�/�/?"?4? F?X?j?|?�?�?�?�?��?�?�?OO0NPO��V@�+?OyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_8�_�_QBDEVYN�P mO�_!o3oEoWoio{o �o�o�o�o�o�o�o�/ASewPALT�q�/x� ���� �2�D�V� h�z�������ԏ�8��
��GRI���� B���j�|������� ğ֟�����0�B� T�f�x�������0�j�R�Z���� �2� D�V�h�z�������¿ Կ���
��.�@�R�ԯPREG�~���� dϲ����������� 0�B�T�f�xߊߜ߮����������X��$A�RG_� D ?	����9���  	]$X�	[M�]M���X�n�,�SBN_�CONFIG �9������C�II_SAVE � X����,�T�CELLSETU�P 9�%  ?OME_IOX�X�%MOV_H����REP�S�&�UTOBACK�����FRwA:\x� Z�,x���'`��xǣ��l�INI�px����l�MESSA�G������A���OD�E_D����#Ox�P2l�PAUSVA�!�9� ((O<������ ��(^L��p��ej@TSK  u����o��UPDT) ��d� ?WSM_CF���8���%�+!G�RP 2
5+ �L�B��A�#�XS�CRD/!15+ �������/�/ �/??(?�����/p? �?�?�?�?�?5?�?Y? O$O6OHOZOlO�?O|(�r�GROUN |S�CUP_NA��8�	r��F_E�D��15+
 ��%-BCKED�T-�O0�%_I_�� ����-r�_x��o�o�x���U2 r_/��_�_�R�o�iUp�_&o�_�_ED3o �_�o�_n_o�o9oKoED4�oro'�onpn�o�oED5^ �:n����ED6��o��npK���%�7�ED7�� ^����n�Z�ɏۏ�ED8J�*_��N_�m����m��ED9�[�ʟm7����#�CR_�����7�ٯD���ū�@�@N�O_DEL�O�BGE_UNUSE�O��DLAL_OUT� ��R�AWD_ABOR�𦾦A�ݰITR_RTNz����NONSi �����CAM_�PARAM 1�9�#
 8
S�ONY XC-5�6 234567w890H ��@���?��( АZ���y�u���\�HR5o�8������R57����Aff��\�L�^� Z��ߔ�o߸��ߥ���  ���$�6��Z�l�a��CE_RIA_I�(%;�F�!�{�x� ��_LaIS$�c%����@�<��F@�GP 1]Ż���O�K�]�o�.�C*  �����C1��9��@Ҧ�G���CP C]���d��l��s��R�������[��m��v��������� +C���& ��G���;�HEנONFI����@G_PRI 1Ż��T� ������ �CHKPAUS�w 1I� ,� BTfx���� ���//,/>/P/�b/t/�/O��x���8�!_MOR���� ��@B�{%���?�̋��	 �"�/:�/.? 9��;P=45�"����-=ֱ?99�D�3�@K�4��<P�������a�- 8��?OO�J
�?KO��'ưS�P1��:O��i]`��PDB� �-�+�)
mc:cpmidbg�Od��C�:�  , ,w����Ep�O-_�C  �  uKP� T�@�Oq_<Z�&Ў&ЏS[_�_V=Y�yDAS[g�_Do�]�,�! UYf�_�KoAMo�JDEF 3ch�)�B:`buf.txtqo��Mro�0����'�	z�A��1=L���j+MC�#�-,���(>ss�$�-�r���Cz  BH3C�s7 C���C��M�F��iDP�E�~�WJ�!0D�tE�q�aEpIJ$��3HHƷ���{G�G���GG���N�[5K~w)L���XWI����du7���4�),�,�.*װ�,�,��@�u��K�x6�q�* ��* e�D�n��pE�WL!0EX�E�Q�EJP F��E�F� G���}F^F E��� FB� H�,- Ge��H�3Y��z�  >�33 �T5�WDn6�P1@��5Y����"��A�1WDq<#�
 �O+�)��Zj�bRSMOFSb���n6��iT1� �DE  �?DR �
�,�;�&�  �@�:��nTESTR�bo�8�R��!�/43�nvC+�A�WJq�E [��rq�C�p)B1 w�Cy�@T�6���T�FPROG %ź��ů���I���𦶠喤KEY_TBL  �6�Q�!� �	
��� !"#$�%&'()*+,�-./01g�:;�<=>?@ABC��`GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?���������LCK�X	���S�TAT*��_AU_TO_DO���G�_�INDT_EN�BK��"R��i�[�Ty2��\STOP����"TRL��LET�E����_SCR�EEN "�_kcsc��U���MMENU 1"~"�  <�� ��|�WE[߅ߺ�V��� ��������,���b� 9�K�q������� �������%�^�5�G� ��k�}��������� ����H1~Ug �������2 	AzQc�� �����./// d/;/M/�/q/�/�/�/ �/�/?�/?N?%?7? ]?�?m??�?�?�?O �?�?OJO!O3O�OWi�;�_MANUAL��Ϟ�DBCO��R�IG�4�DBNUIM�`�<q*�
�A�PXWORK 1#"�ޟ+_=_L�^_�p_�[�ATB_�� �$"��ipT�A_�AWAY�C
�G�CP *�=���V_CAL�@M��R�BY��h�*��H_�` 1����� , 
^@7�6�Boo�f�PM���Ij��\@��cON�TIM��*�ɼ�fi
�$cMO�TNEND�#dR�ECORD 1+�"�er9�Q�O� Oq=6��R{��� Hx��O�s(�:� L���������ʏ ܏� ���$���H��� l�~������Ɵ5�� Y�� �2�D���h�ן ������¯ԯ�U�
� y����R�d�v����� �����?�����*� ��N�9�Gτϧ`�^�� ����=�������(ߗ� ��^�p��ϔ����� 9�K� ���!�H�� l����ߢ��K�a��� Y��}��D�V�h����RTOLEREN�C�TB�b�PL����@CS_CFG� ,0k�gd�MC:\��L%0?4d.CSVi��P�c���cA CH
 z�Poo�n"W�^m�c��RC_OU/T -�[=`�o~��SGN .�U�r��#�2�5-MAY-20? 15:37 �Q��
1:00 af? P�X���n �pa�m�?�PJP�{�VERSION ��
V2.�0.11�kEFLOGIC 1/�[/ 	tH�P���P��PROG_�ENB�_r�UL�S�g �V�_WRSTJN�`�Fr��TEMO_OPT?_SL ?	�Uac�
 	R57Y5�cO 74T)6U(�7U'50y(t"2�U$tH�/z2$TO � >-�/{V_V�`EX�Gdu3PATH A�
�A\�/]?o?�kIkCT	aF�P00g��Tdceg���1STBF_TTS�h�I�3U�Cda:�6�@MAU �.�bMSW��10i�Q<�l� ��2�Z!� mO|3bO�O�O�O�O�O��O_tSBL_FAUL� 3�_�cQ�GPMSK��bTDIA��4�=�d`���a1234567890�Wc|6P�/�_�_�_�_ o#o5oGoYoko}o�o��o�o�o�o�o\SpPf_ *��OR*� ?%�PBhz��� ����
��.�@��R�d�v�H|��UMP�4!Y )^��TRpNBKS��ĀPME�5~ЏY_TEMP��È�3��D3�����UNI.��YN_?BRK 5�����EMGDI_ST�A%�W�NC2_�SCR 6G� �_����͟ߟ�f�����0�B���~�e�17 ��;������¯,R|�:d�8G��a� ������N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� 0������@$<��)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� ����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/��/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgO�/ �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo�Oqo�o�o�o�o �o�o�o%7I [m����� ���!�[oE�W�i� {�������ÏՏ��� ��/�A�S�e�w���𛟭���קETMO�DE 197�.v� '�� ��W�RROR_PR�OG %�%����X�'�TABLE  �A��������њRRSEV_�NUM ��  ����)�_�AUTO_ENB�  #��j�_N�O� :�
���  *�F��JF��F��F���+E�p_�q����HIS��h���_ALM �1;� ���F�F�+�� ��$ϐ6�H�Zψ�_�%�  �D����ې�TCP_VER �!�!F�j�$E�XTLOG_RE�Q������SI�Z����TOL  �h�Dz���A= ��_BWD�5и�a�	�_DIO� <7��	�h�<�k�STEPw߉�|ې��OP_DO���4�(�FACTO�RY_TUN��d���EATURE �=7�a���Handlin�gTool 7� �DER En�glish Di�ctionary�=�7 (RA�A VisS� M�aster0�>��
TEa�nalo�g I/O7�>�p�1
a�uto �Software Update��� "`��mati�c Backup~;�d
!���ground E�dits�  25�LCame�ra��F�� "L�o��ell��>�Lw, P��ommj��sh�8�h600�%�co����uct�%���pane6� �DIFD�'�tyl�e selectv�- `�Con��~j�onitor<��B�H��tr5�Re�liab�� �(R�-Diagn�os���:�y�Du�al Check� Safety �UIF��Enha�nced Rob� Serv��q �(V�Use�r Fr���T_�iE�xt. DI[O ��fi�� Z��\=end Er�r��L��  pr$�[r��C  P����ENFCTN_ Menu��v�����.fd� TP �Inp�fac� � 
v�G��pl�k/ Exc	 g5t����High-Sp�e Ski��  �Par\�H��G m�munic��on�s��\apur�� p���t\h8y��conn���2� !D�Incr� strZ�i�<��M-6< KARE�L Cmd. L�� ua���8sR�un-Ti4 En�v=�(mqz m�+���s��S/W=�"�y�Licen3se��' a����ogBook(S�yo�m):��"�MACROs,~�/Offse��f���HG R��M�1?�MechStop Prot���d 5
$�Mi�eShif��9�B;6SD�Mix �����7�y�Mode �Switch��M�o����.& �MT�&��g' 65�?ulti-T� �����Z�Pos��Re�gio�  ! �7Pr�t Fun<b>�6iB/1���Num ��dx�P�`�312  Adju<:�/2HSM7Z*� oY�i8tatu�1<�AD RD�MotN�scoveW� #��3��uest 867.�9oG � �?SNPX b���<�Z#LibrV�;�Ort IE,� S$�@�.�0�� �s� in VCCM,9��0�� ��!�9�3��/I� 7�10< TMILI�B�MJ0,@� �Ac�c����C/2@�T�PTX"+QTel�n �Lq3�%|(P�CUnexc�ept motn��� �0�0,	7�\m72f�+4�|f�K  h64aVSP CSXC9���@(P�U["3� RI�N�We'50�,D��Rvr�	mcenS@� �QiP^ �a0��3fGri�d�1play F� O`�fp@��vVM�-�@A(B201� f`2� ORD�|�scii��lo[ad3�41%�lJ�i�Guar�dP�m�P��k7�b]aP�at�& 0N"Cyqc��0ori����`iC00Data�@qug�c�3[,�`�3FRLOAam��5<�3HMI D�e�2(�1oc644��0PC�sePas�swo�aA)qp�1pp���{-+PvenjC�T���YELL�OW BO�I t�"ArcV0vis���%���Weld�� cial�$  �  �et�Op�A ;�41\\�5a 52��a��po)@`@L�aT1���50.23HT� @ xy�R:�#82���`g�P���xp�� 12�AJP�N ARCPSUg PR\A�TEh0�OLwpSupg�fil5p�Q��^ l�wcro�6 "T�`Ч3ELdx�!��SS�wpeetex^$ [J3�QSo�t� ossag�% T��eBP� ] !9M�ViCrt��39�V h	`�stdpn6��r�o� SHAD�pM�OVE TF MO�S O � D�get_var ?fails ��ߐ#  � D��E���� Hold Bu�stdCVIS U�PDATE IR���CHMA 62|�q�WELDT�@�S ) "���:� R741-�ou�
�b��m BA�CKGROUND� EDIT Ò �m41�0REPT�CD CAN C�RASH FRV�RTO�Cra.�so 2-D��r �0�r$FNO �NOT RE��R�ED � PCV�l�JO�P QUI�CK�OP FL�EN .pc�c����TIMQV3 �ldm�PFPLNs: 燹 pl 2����FMD DEV�ICE ASSE�RT WIT i�C��sANġACCESS M �uaŀo1Qui��t<!�C"�USBU@�- t & rem�ov��<�2� SMB NULApܡ���FIXW��HIN�͑OL2�MO O�PTt�PPOST4wp��D��- � �7Add��ad. 	�[io��$P:�Wu`k.$ѠO��IN���M��CP:fix� CPMO-046 issue�t�JСO-|�2�13�0���SET V�ARIABLESxΐ�$O�3D m�"?view da`P�Wea�80b. o_f FD ��u)�~�x OS-1�p� h s v�D�5�t��s ��lo ��(� WAx��"3 CNT0 T�fS$Im�Z#ca���PSPOT:Wh��p��s�STY܄A�t�pt�do �GET_l���VM�GR LO�0RE%A�pC��M`P��@ Y��0�ELEC�T��L��ING �IMPR N���R�ɰ̐sPROGR�AM�RIPE:�STARTU�@A�IN-��D��QAS�CII�d�OF �L���!`PPTTB�: N��MLKdmie�4��:�moW�gall��R� Nu�:Qr� Ang��郲`d��tho�n[� ch >`ܐ��r R2toun�H8}5@�iRCalA��"Sign�0�pI�,A�Thresh�123�#.c�H�ڰ : MSG_9P�єper �ࠡz��A�zero5P�� A�  J�!O�I�mr � 2D�0rc� imm�`SOME�s�ON�����>�0SREG:�^�5� LB A9�KoANJIH�no��r�`c	��n dq��� -1o��IN�ISITALIZ�ATI��weX��0= dr\  f���aP���minim�90rec 1lcz0�:?!blem��Cro��L�<3a iң 09 ��b�d�w�-� ݡ�0�w ulHQm@se�4SY��M��s���QЧ 09�0�Wlu� E;BR%e��jձ4�1���3m ���Par�r@ �G�Box fo �TME�ːRWR�I<���SY��\kڼ�F/�up��de_-rela2Qd�|�#5�betwe�p�IND��GigE� snap�us�5�spo V�T�PD��DOs�ġHANDL �`�Q��i�D��n�0 f.�v���Boper�abil�` tm�CQ��: H5@�`l��L�
! ���m@ph�s UIF6L�PO>�FA�����ΑV7.��CGT��pi�AsM�5pj��)@U��ine-R�emarkO@0 �RM-�$ÔPAT�H SA̐LOOqS���v�`fig�GLA  �0%����p��J� ki q�t�her�A� Tr�`in�DW����2�7�� X�е����8`n;� C� ��:�  6�d� y* it� 35\k�Pa�y�a[2]_�D1�: g�s> do9wD2	SDISp�1��EMCHK EX�CE ֠�$MF I+  ��h�"�P�4�Վ�B0 ce1�Ȣ��me�� �c�� !?��bP�� B�UG��yB
�@DŠPET��V0�0�T�93X�XPANS�I)�DIG��O�  H5�P�CC�RG ENCCE�MENT`�Mm�K� 1A�H GUNOCHG OA�1Tڐ(����Sg\d����10ORYLEA�K������LC �WRDN R��O�`j5`PO�SPE�ްCG�V ont��VM����W��.@`GRI,@A�7���� �PMC ET�H�0i�SUذ>� �H57�P0PEN�S!�N���ː RwE (i�ROW<��³RMV ADD�  II�=p��DC�^ q�T3 ALA�Ӏ ��m��VGN? EARLY>���f n� ��衸E�AL#AY7u�СPDg�ˀ�H1SS8�OUCH��D��Fh�����P�CDERROR*PD�E��� WRO��C�URS�PٰIp@N� gҰ�?Q-15�8Kwa���SR ��ġU3��\ap(tp��@T�RF@�R �\`�UB�U �`���#RB�0SY RU3NN���`10�ఱ�BRKCT@qRO`q�Ԁ���CDAX�x�Djj�EISSUcpހ\��D��TSI�a�K�tXM�IPSA�FETY CDE?CK "M6��� dѤ�[`S U�)��4}P�@QTWD��E�'QI{NV��D ZO��ࠂa�sb_aBDUA�L@|�'QòF��EԨ4l�6��P`NDEX F�P�U���SUF�rPk�Lbѳ�R�RVO117 A�y�T��챤 ��FA}L�BTP247��r�P?q�EHIG�P�CC n��0�ESN[PX*PMM�Q ��)!SQ�"V��8T�b|DC�BDETEC��cds!Sˀ�BRU/b�63���s� 02"��t�s�'�!h� Z�T�7pS��"e���߆��,����߉ـ�0��
ա��ق�csc�r�ـ �dctrld.؁���fIّ��!���fـ\*��878��-�%� ��� rm��
��Q�R��78�RaIـA�̑ (���~��Q.����ao�ـ\ ��a:P���a��I��=ta 3 "K:���a�<�#�o��tp؁ "PLCF"E!x�ـ�plcf��p�ـ-���mai�ـN���ovc���ـt�/�ـ�������ޢ�r674��Shape GenwـI��R,���ـ1T�іV� (5�ـ��II���� �+��Xـl���sga 4Pg� 4j�I�r6ـ�Ų5=�5ѺI���e[ts6� " PC����nga�GCRE�ѿ|�5��@�DAT0j���5ŝ�t.!���5�a񯜳A�gtp�adb���Y�tput������ñ�ց2ـ��5Ĺ�����s�l�q� 7�he�xy��4�����2�kceyy�ـ"�pm�������us9ߜ�gc ـ����+�H��a�j921��pl.Colly󔱾��r�ВN��ڕr� ({�ـip���r��('���8�7=�7����tp�� "TCL�Sj�|���clsk誨D���s�kck ���)�U������r��H���71a�- K�AREL Use� Sp�PFCTN�j��7��a�a��� (��ѡ�� �ـ������6�8=�8"  � �ـ 0S��(V�  g lm� 6�99��~ F�)vmcclmf�CLMl��`���60vet���LM�:����sp]��mc_mot���`ـy���suX���60���jo�iT�J��_loqgH��trc��ve%�� ������g�finde�r��Center� Fb!��M�520�����g��  (m)r1,���fi��1 ��a#z�� �ـJ���$tq� "FN�DR����$etgwuid@�UID� ـ
?1��E7�q1nufl�6 �ـ>_z#ѯ7A��x��(�2#���$fn�dr����c$��tcypS$]�CP M� :H�3ـ517��g�38�vC�gD�* Y=�F| Ց� ^ ��&�CtmgA4�P��O �CG1ՑO7�Y��8��Etm �?�Wـe0�?�C�Rex�ے����Z��ڔXprm�؁�_�D�_vars�_Z$M���Vh@��0��`�gG��ma�w��Group�@sk� Exchang�{@ـÖMASK �H5�H593 MHa�H5���`6�`+58�a9�a8�B�a%4q2���b(�o�#
k�/�غ`hp8�0�Y0/_цt�qTASAKY_�r��pz�h��Z�m@��������SD�isplayIm���v{Gـʑ8�OJq(P%���@a���a�� ـlq�vl "DQVL�t���q�����Ϧ��y�����1avrdqq֏4ᩅsim����0��st��o��d ���������v�0Z�𨁯��"v�Easy� Normal Util(in4��|+11 J553��a�c���(���0���)�M�<�O�<� k986TA8��#�4�� "NOR�
��1�_���|�su��.�������7���a!g�y! �menuu��g#Mx�����R577� �90 ̒J989F��49�L�A0�(�ity�E�A�,�P�m&��mh8��"8@ 2��܄����C8_�Sշ�n "MHMN�r%.Ը%���ͯ��s����i�Ը-at �Х_�������ֶ��#tm�?мz�1����"Q�2�Ͽ�z�3zos��odst��
�mnx�O��ensu�	Lm���hRaL�߃�~�huserp�a����c~���Ը5��ɯ�����oper����XԸdetbo `Ý~ ��LUA���������dspw�eb���+�X���u<1��101W�הּb�2N�A�e�30A#�0����4N�;2e�5���|����"��CalxN�0�O��Z��0�O��$�S%j{�u���? 0S�}����ump��\bbk7968�!68�!���b�eq969�9��%��F0b�� "�BBOX�ۍ�s�ched����s�etu~Xk��� ffH)�0�eq)8��0�col(�1�bxc��8�li �Љ�aI���W!i��e@m�rof$TP �EB!TA&@ry|M4127�*l!(T\�Q!RecX"H
�qz�?$�it%�?#сk97�1�!71�{�F�$p?arecjo��A���?'����Xra{il�@nage��~@]��D2E� [0 !(?:H͒V|x@1ipPMa���3�p�!4�"�4�u��3paxrmr "XRM$��3�rf�Ͼß1��1ꫝ0�yturb�sp'G#��^@ �0s15: ��625t/ ~A��\BH�'ZDiy!:k�E�6�"A���H� �7��P�.�E!�pd "TSPDx�}�T�GtsglD���kY��O�CiCsRc1t%���HvrvQ����K�P,��A  �q#-a21��Y@AAVM� �r-b0 �fd�E`TUP him� (J545� l) �i`616� V2VCAM� .CLIO] Y10k 5W`� (F�`MSC ����bPs�STsYL�Sua28 kr��`NRE I��`S�CHgRpDC�SU tpsh ORSR ��ua04�EI�OCW`\fx�`542 LEX"�`ESET��iay`0�shi`7y`"ROMASK�b7o�.-`OCO[�x�a7p�3Sv q`t7p0kv6�U`xv39_v�xLC�HRvOPLG�w0=3;uMHCR3Mp�C�`YaP`�p6�.�fia54; #�MpD;SW�`588�ip�1�a37 88 K(Dr0c�5r4��N�r7 qj5r5��5r^v�p5�"9�PRST VR/FRDMC�S�a���-`930 ��`N�BA  g1�`HL�B 3 (�aSM޹� Con�`SPgVC Lia20�#�-`TCP ara�m\TMIL� r�PACC�T�PTX �p�`T?ELN 96�0�r�9/uUECK�1r��`UFRM et�L�aOR ���`I{PLKeCSXC�p�j�qCVVF l� F7�HTTP �strbZ0zcpCG�y�8�AIGU�I�p7 ��PGS �Tool�`H863 dj��qM�Ozq3
vJ684c�\$���sق�s'��1ےs�a96 TwFADȑ651�Cnq53 � oo�b�1�44r-�k�r9��VAT��J77�5 �R�6uAW�SMے�`CTOP1 �q�`old��a�80;!diy�XY�Y�0 e��i`8'85 '��`L�`u"Խ`� 7H�`LC�MKP��pTSS �J%�
�W�CPE� \dis�`FVgRC m��NL��U002 
�en�%�6 65Jr'�7[�U0�po�ࠠK�2��t� I�4 URI��5�&�U022 �nse�{�3 A�PFI�`{�4�2��`-���alOP��1�C�33O�͐tpt�sD`U040g�4�3�ٲ4�۰j� �"sw%�1`b	�4��C	�5 ��wx�5=7�eU061��S�]6ұrob9�5g�i��68����!!��	7�w�7�Ё�%���_"rkey��3w���4?ǽ���T���8�'�089�U09Ȯ��P��9:���2 �&�l �9&�l��9�B�VrU15�P�M� slA �3#�}�R��1q�0v4�7��/108 	�eэp�hc ��s�1�q�4�+�1����A�5/�tRx�1����1]pu�Qѡ�t�1�����`��)3����6��1!p ��`�о�- W8�1�47 ase C��U`sB�1 82���1�4�8 (wWai��59 �N�aU166�W�1�"W�4� j U�6�#U�	7�3U�8�3ѱ��B��1{��2 ac�t���6 "MCR@�ِ4�1�������967ǑU193�3��6��2Y�sP��2A��21��as� F���<�2-���NE�2 wF���55�T(��� ��cر5)��w���q��p����qf ��L��$������q4dB��2g�8q��8�51��""]�}�q��< b������B]�� �f�; `�̑ � 8 16 (ݰ�BA ��AAҰ�]����g :�!��`8 bbfo=� t� j�� 7 \� ]��� �2 k_;kv��74 &!�����W0H5��57>&�579 h� L82 %"���4 3��5����5���1��594 �U219 7,-�6��p��6i�\tch�H6ur% �4S3� 90� h�&>�\j670��q���r!tD�4�h�&�t�sg��lc�S�FrE�H���#F�����hk$�� sC�� ���"F�L��df�lr��� �� ����fu!l%�gvPva����sA� ���"D��3��!creex���!�%��!�%�,���6j6z�s�!prs.�! �%�!5�hA�P 5�fsgn��/�/�,at<D�AD����qs`R svsch�`@Q!Servo �S�!uleoCA5SVS�!44���F̝�1 (�0Ached�0,1�EA���� �2Q��0��^��r0�U)1BBc��� 
%P5)Q1�V-#�3��1css "ACS�WVY88"gA�`8!�/�0��@e�Ҿ#M���C�3�torch�m�0�- TQM�a�1�1M%'�9 J�5lA598 א1
�!7)P8<P(1̢A��ء%R1Qte,��!)E A5E`ASv��s mLC6ARC_�� 1�4q� X�V�Ht!tc�A�p�Q�4��R F1j 7T!2�SEPBpPQf-!�RtmkQ!�p@60X��/�PRC 8S�Q#�S�) P�2a�96xAn`X�D.<bH5�1�U�}E� T�Qf#` aQ!<���F!�T�!!�a4�3FcRO�Ttm�R!av`58�_�WP��MA$q�E8��>rp�in_���o
�@e`AcB�rr�)u8�!�U�etd�ѧ|�U�Qoveto�#�$,�S�mmoni�tr42�=�Q�c�st,"M_va�P47M��V�0�! 5�q����ameQ!Ɂro�l�A��43$Q0a  Sp��1�01$P�25�AKR  ��� 0S�(V�Ɂ)xj818\nl`mD��zN��r>�MPTP"�O�>�qmocol�]/ 
�Y1�4Xa�@��2�0�i�53(1��Touch�!sؠ�2%qD2J5 !IU�٠��= b�0n��A��]�vP����z�EOWJ�th���Kwc���{�e�tth8!THSR�Xâm�t�o "PGIOsRd�'z�;wk� "WK1�avL&MH�PH54�%5�Q5�o��m`A��Bq@7z@6���18�ap�PMor��tsn�@T�A�o�c���"�����m�uA��T��p���T?�|�$m4�TM�!2�54�>� ���m9�w�f��S�3G�qor�3���"641���8ⱐQ!A�,HE!pRU <��m�Re�h-g "�SVGN_��(co?py "COTA���U(��r#j0 "FS�G��_�eh��f�@wA�SWwjRbY=sgatu���!��;B�tp�ATPD47��9 a79s��̠�sg8!��GA�T&o<Rc9  �Ħ�1�t2`%1�&��1�bpv�1� �&�1��B �1� 6�1�chr��1�|v�1�sm��1�v���?gtdmenps1��(v0!1��mkpd�t�r1��]A1��pd��1�$&�1��mvbkup.1���6�A��mkun̠�G�pr���mk�l1�e�P�s1�nix��0&1�ldvr����glg�t�1��&����#�auth�.p�&��1�����) sud�1�7� 1��G�1��\1�g b2�p�w 1�6O�Ł4� 1�Ђ   946"1�����1�t\pai�c\p4k947�1�wc��1�icgtas-�Mpa�cck0m	�	Ngen!1� �wl��Q� sctfq��q�wb�����������vri/�4�^��B1x�D��Pflow�@6��Ac0ow�3<R50?���Q�TR�  (A0e T�)B�Ԗ�cud!�w�1���z�ac�$046` a� =�f�+pa`Ra���!1�355Ţ 1�F�ѡ�)a%��;:�afcald� @�&�0����%�f�m:�"�#�4�`��'a`"�3U���$�B1�! track����@aine/Rail TrP��{(s69�/�@ (L ! iEYB�ʔ_VB!BHu��a YB38P�48'7�	�F2��4���/�C�B1�3Ţ3��/�IUal��1�N�T����VA��zQinp�p�?0HVaen0 �?DXWApuA�YqBzQtstd�0U�@1 GW ��]�j�VD����E&��VH@���ope/ners^CO�`�AGDev/w'~6�F�8��񭁶��bA�aes�#1�]�ג�d�`���m�d1�k9�@
7�6��#1��/b�e�paop`aOPN��Wj�`��Krcel}?�Exg���Y`5Dv��tscx?t��a��s Fuvrop /�Dw�nDh��b Ar5��QB�g�dk�j!>�� Pumpv$A� ���/�1�a;��M��T�q�i���t��4U�1� 0S���O \mhplug�gr7Gh���u|bZ#��ioh#Cp{p��v(�ALIO1�51�@7��93�QE51�91�����4��� ST�
R�t�J�989��/RLSE(�g1�@Cd�(M�1�/O�'�Q�)�D��G�1 zq�H155�'?��zq�tcmio��MIO�$��tc�q"CL01d�UQcP�|�io��u~0%�l9�zp���v�1o���Q�tzt����dtz5I$���V%�rh#Inte\�Q�� Co~Po�q�vRP1�hd�B55G4 (l�oBv�,�Q8�H��Tcipc�oo�&ڱp5�A�(
��������"7`���5aڰd�QCD�W�	�����8��ڱ�rcnQd�_׳1p�a��ײ������S��a��O�2kz�rpcrt�ᱯ�pٱdEc��S d�\����u�E!߳vr2k �pE A�-�x�_B\"� gchoO�l"uC��8Y 1খ630@ᗷ �@�� �ӿ�q��ԑ��GTX�? �Е1chp "��XOh:�3�&�"5x!E��\p3 ���P��j��d 11�$h��Plao���ұ�ch��3��s1��a��01���#Ar��0� !oCB��spq[Jm:�k�7�)�vr�Ҿ���pa!X%-J�FRAJ�wWatpqrnev' �����fQ��D5�`��.KrboT ,�$��PG�[!�sm�ICSP\QQP5y��!QP����j�H51z�9%3QP7y�6����d����5��R6QPl���NPR�`(P@a/am S`u�b��|ĉa4tpprg�p��B�	�Z�qratk932(q v��/sc "iC��~�atpr�_�qq�z�;F�LGdsbl�flt{�ёsab?le Fau`���CPav�aQ��`aD�SB (Dt$�t �d�A����QPh"�E1��`f$*��3[S� A6�"tdj  "PaV�Ohf$�1sbj!��1�"\:1gc��.�f%�d�u�550^CAdj�ust Poin	t�b��J/��-�0� �4�a昐A��j�O�N/0\sg�4��wު1\ada��"A�DJ�M�j0�et�sham�SHAP80���XDjpo �e� �G�a��UGQPG'.��1�:�k@ab5�J�KA�R`�iagnos�ti��!�a��66C J�C��a=P(Q�L�Q&T�o�fkrldeP@���	 ��SHQ��)�3/ρ[pp���DBG2t�!O ��U�Rѯ#��V��F( `�шS7��Q�ip{��M�ipper �Op��Pq����78? (MH Gw�1R lbk_�fTcBQ��0&,�d038<B8t��(E��c�9_9t��$Tc��k����8$q� SdrnpVǁ��Qd��Ő6Tea�=���r �Mat.Hand�lv �an`W�� M�PLGv�A_�p�q( �sє�f����g�� b��a���f���� ��>@$w����Dw��@EI d���uu�m����fhnd "F~��  ���
��#� ��p��>��7(Pa�0To@�$V(�!!�3#p��a>���{�Q�k925��2�6�q�3�{�p����2p	ş�y���gse>0�GS�qďėPR��T`���a���tp��<��{�dmon_�q��Ŗ�ans���vr ��{�=�����ͪ�<y�֯wsl� � pen��D��Y�WA��823X�Q
�G�0! '�&P��8QqIQ�G:Q �\sl��!q ��v���������֐��_�`����"SED�GiOٳaQ�tdg�@T�AF8�F���BN� ��ÑQm�7���ڱA��g;Ж�Q�����q�NS�ileg�y�e�� �ϟ�9�F'QQ�LaQQj517So�3-[�JV�?�'�#4A�49GA�WL�aw {��no�Qfԫo�H17@D�#a�����0t�?  >���LANG j�A5��5�5� gad5��C5�TC5�jp .5�ce���5�ib=�5��#5��уpa5��C5�WҸ�j�539.f5�]QR�u5� Env
 5�5S��K�3y ��J9$5�.� �;(��G5�2D25�JS���p(K}�n-T�im��"���"��3pH􅓹���\kl5�UTIL"�����?r "QMG��,qp5�C5��1 "5��ړ5�s5�\kcm�n��+��r5���u�tM�_�lread���ex����"��E\��l$"��135��rt[! -5�tu@va��`_��5� �`cCV����\p ����Bp9tbo�x��_qcycs�}kRBTvve�riOPTN v��l��e���K���hg/�a�gp.v1$�"1$p�tlitDP�ND�BPm$dn#te\cym$8$o"��#mnu3�/�/�/��.5�/�/m$��UPDT ite��>.3 swto95]�-4oolBD5wb95���-4FR-4Y�� /2grd�-4��-4�b-4��w-4B-4.3��-4��-4'�-4�.3B0l<� /2bx "�5�Q5I.3tl�7��AE�#/2r l\�6�@Op�-4 :4ColD5eMa-4+�C�5K�-4�W�Q5ml�-4Cha�ng95}�95�qQ5r�cmdE�b�OZ�`6 �5,r�7�6��7�5&rL_+]22=_O]2� �c_u_3U4<_N^57x�_�_1UCCFM�E|y��_accdau59#�6cAEX`�/2|@�Da��4|aO/Jm�a �5�-4@�4�aAOSJ 	Q�e�o�oY��`-4��ZDQ-4sk��?�@rtet�q-4\$x�3�q�eunc.-4p��4�q�5sub�5p��5E�q�5cce� @oRf^opm4E�o�fv�7�o�eT �c�o�n@t$
Pte;�q �@��f\��k��6;�-4/Ѓ -4K�D�x�zh!-4xmov�b�q�et���f�"��tgeobdt.8���ƥ�etu� ɐH��ɐ��tɐٓxߟr�z��var'���xy&��pclBJ�cɐ��ɐ�eɐ?gripsu�����uti�����in�fpo��ܯ�ɐ������\����ɐ(�Ʊ�8�p��n��ɐ%�ɐZ�mT���ɐԶ��\�ogġ�Ʊ�%�p�\�palp�����s����ɐݵ��Ŵ��⩚p�p����pka�gd�%�7�lclaAyY�k�A�ɐ��dɐ5�p�������B�� |�|�������q�����rdmͿ��rinT�-�?�sO�Q�c�̿b޼s���ߧ�tv����h���stn([`��tX01ɐ)�aDɐ� �Tul4��q��g�26Ϥ�up1d����vr����נ1}�3�נ��ϵ�gil3C�U�l4����T�5e�w�s ߘ�8֠�߻�wcm�(��xferϪ�t�lk2pp��c�onv�朗cnvݑ��5�ag, y�Glct���n�p��nit0���d�x��(��  �ɐ� 0S�(V��U9al �pm�Wse��2�� ��V�C��(�z���A�0�|�m����&$��޷'#ro��T/f(&���p1�mI��, ��$�+���/�)G��?�+�� �L�ɰm  ∡P?b6D�4rg� �����������? �9�� O�7���� ��>�/�T�a�8/ �C�����E��b,֡)?�*��nq?_9l��-!H��  �>HA |�p�QU?1 p! O���v�P ��S 	�QڗR@t�`  �?��ɐ8� �M<�.Oreg.ԃnO~�o99 ��� ���$FE�AT_INDEX�  �S ����P�5`IL�ECOMP >����ba�Pa�RUcSETU�P2 ?be~lb�  N �a�Uc_AP2BCK� 1@bi  �)�R�o�o  %�o�o�Pe`�o)oe �oU�oy��> �b�	��-��Q� c���������L�� p�����;�ʏ_�� ����$���H�ݟ�~� ���7�I�؟m�����  ���ǯV��z��!� ��E�ԯi�{�
���.� ÿտd�����Ϭ�*� S��w�ϛϭ�<��� `���ߖ�+ߺ�O�a� �υ�ߩ�8߶���n� ��'�9���]��߁� ��"��F�����|�� ��5���B�k����� ����T���x��� C��gy�,��P��qi�`P�o� 2�`*.VR�H� *Kq�0w��2PC��>� FR6:���/�T@`@/R/��=/|,C`/�/�G*.F5�/�	���/ <�/$?�+STM D2M?X.�E?�=�� iPend�ant Pane	l�?�+Hz?�?j7�?p�??-O�*GIF7O�aOl5MO
OO�O�*JPG�O�Ol5�O�O�O�5_�
ARGNA�ME.DT?_�"o0\S__� �T�_�@_	PANEL1�_�_%o0�_o�?�?�_2orog`oo/o�o�Z3�o�og�o�o�oH�Z4zg�h%7�KUTPEINS.XML��o_:\���qCu�stom Too�lbar(��PASSWORD�~�FRS:\k��*� %Pass�word Config�������� +��O�ޏs������ 8�͟ߟn����'��� ȟ]�쟁��z���F� ۯj������5�įY� k��������B�T�� x�Ϝ��C�ҿg��� �ϝ�,���P����φ� ߪ�?�����u�ߙ� (ߒ���^��߂��)� ��M���q����6� ��Z�l����%���� [���������D��� h�����3��W�� ����@��v �/A�e�� �*�N�r�/ �=/�6/s//�/&/ �/�/\/�/�/?'?�/ K?�/o?�/?�?4?�? X?�?�?�?#O�?GOYO �?}OO�O�OBO�OfO �O�O�O1_�OU_�ON_ �__�_>_�_�_t_	o �_-o?o�_co�_�oo (o�oLo�opo�o�o ;�o_q �$� �Z�~���I� �m��f���2�ǏV� �����!���E�W�� {�
���.�@�՟d��� ���/���S��w�������<�ѯ�Ơ�$�FILE_DGB�CK 1@���ʠ��� ( �)
SU�MMARY.DG<篓�MD:�[����Diag Summary\��i�
CONSLO�GQ�4�F���߿n��Console �log�h�G�MEMCHECKտ輿J�c��Mem�ory Data|d�l�� {)O�HADOWY�>�P����t�Shado�w Change�s��£-��)	FTPҿ?���C��n���mment� TBDl�l�0<��)ETHERNETaߑ�"������n�Ethern�et ��figu?ration��s�~V�DCSVRF`�pF�X�q�t�%6�� verify �allt�£1p=�1�DIFFi�O�a���u�%��d�iff���"�6�1p������{� ������	9�CHGADE�W�i���u��&��9�2�������� �����GD M_qu�.9FY3����� ���GD Ugy/u�6/��UPDATE�S.U ;/��FR�S:\S/�-o�U�pdates L�ist�/��PSRBWLD.CM�/�"�/�/��PS�_ROBOWEL ��g�\?n?���?���? �?W?�?{?O�?	OFO �?jO�?{O�O/O�OSO �O�O�O_�OB_T_�O x__�_+_�_�_a_�_ �_o,o�_Po�_to�o o�o9o�o�ooo�o (�o!^�o�� �G�k ���6� �Z�l�������C� ���y�����D�ӏ h�������-�Q�� �������@�ϟ9�v� ���)���Я_����� �*���N�ݯr���� ��7�̿[�ſϑ�&� ��7�\�뿀�Ϥ϶� E���i���ߟ�4��� X���Qߎ�߲�A��� ��w���0�B���f� �ߊ��+���O���s� �����>���O�t��������$FILE�_ PR� �����������MDONLY� 1@���� 
 �5�Y�0}� =f/����O �s�>�b t�'�K�� �/�:/L/�p/� �/�/5/�/Y/�/ ?�/ $?�/H?�/U?~??�? 1?�?�?g?�?�? O2O �?VO�?zO�OO�O?O��OcO�O
_��VIS�BCK������*�.VD_[_�@F�R:\F_�^�@�Vision V?D file�_�O �_�_�Oo�O)o�_:o _o�_�oo�o�oHo�o lo�o�o7�o[m (� �D��z ��3�E��i���� �.�ÏR������� ��A�ЏR�w����*� ��џ`�����������O���MR_GRPw 1A��L4��C4  B�9�	� �񝯯�����*u���R�HB ��2 ���� ��� ���ݥ��������� ި%�ߤA�5���_�J��Kw��I���Hv��T���^R�<�Q
��aM���q� F��PH\
F��{�;���;U�1�@/�~��@��S���S��E�� F@ %��5U1ŝ�J���NJk�H9��Hu��F!�_�IP�s��?@��u�ÿ9�<9��896C�'6<,6\�b���B��$C�rC��C�2�&B�M`C�&����A�7��Bk�B|���A�v�B+
kB<���������9�A�?�M��r����߁ߺߥ�O����AG�q@5� �߯����4��X�C� h��y��������v��BH9� ��8������{����F��X�5�
��P�X�P�~�`�w������B�����M�@�3�3��������U�UU!U<�	>u?.�?!����k����=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7�:��7p��D�@ ?D�� C�@�U-C��CΏ�'�� �����-�/�C/� #/1��/Y�/�/�/�/ �/�/�/0??T???x? c?�?�?�?�?�?�?�? OO>O)ObOMO��N� P�^O�OZO�O�O_�O +__(_a_L_�_p_�_ �_�_�_�_o�_'oo KoXi�Xo~o�o�oi� �o�o=o�o�oB T;xc���� �����>�)�b� M���q���������ˏ ���7�/{/%/7/ ��[/��/ܟ�� �� $��H�3�X�~�i��� ��Ư���կ���� D�/�h�S���w����� �O㿩�
ϥ�.��R� =�v�a�sϬϗ��ϻ� ������(�N�9�r� ]ߖ�]o�������߷o �{�$�J�5�n�U�� y������������ 4��D�j�U���y��� ������������0 T�-��Q��u��� ���ϟ5GP; t_������ �//:/%/^/I/�/ m//�/�/�/�/ ?ǿ !?�?Z?E?~?i?�? �?�?�?�?�?�? OO DO/OhOSO�OwO�O�O �O�O��
__._@_� d_�O�_s_�_�_�_�_ �_o�_o<o'o`oKo �ooo�o�o�o�o�o �o&J5nYk �k}����� 1��U����y��� ď���ӏ���0�� @�f�Q���u�����ҟ ������,��P�? q�;?��[���ί��� ݯ��:�%�^�I�[� �������ܿǿ �� �6��OZ�l�~�E_O� ������������2� �V�A�z�e�w߰ߛ� �߿�������,�R� =�v�a������� ���'�I�K��7� 9�?���o������� ����8#\G�k �������" F1jUg�g� �����/�/B/ -/f/Q/�/u/�/�/�/ �/�/?�/,??P?;? t?�?MϪ?�?�?���? Ok?(OOLO3O\O�O iO�O�O�O�O�O�O�O $__H_3_l_W_�_{_ �_�_�_�_�_o�_2o Do�eo/����oe��o ���o��
%o.R =vas���� ����(�N�9�r� ]���������ޏɏ� �׏8�ӏ\�G���k� ������ڟş���"� �F�1�C�|�g����� į�?ԯ�����?B� ��;�x�c�������ҿ �������>�)�b� M�_Ϙσϼϧ����� ����:�%�^�I߂� Io[o��o�ߣo�o� �o3��oZ�u�~�i�� ����������� �� D�/�h�S���w����� ������
��.��� �'�s���� ��*N9r ]������� /ۯ8/J/\/n/5��/ ��/�/�/�/�/?�/  ?F?1?j?U?�?y?�? �?�?�?�?O�?0OO TO?OxOcO�O�O�O�O����$FNO �����A�
F0Q� P T�1 D�|���@RM_CHKTYP  �@�����@��@��QOMP_MIN�"P����NP� � X�@SSB_�CFG B�E? ��{_���rS�_�_�ETP_�DEF_OW  ���-R�XIRC�OM!P�_�$GE�NOVRD_DO�CV���lTHR�CV dedd_E�NB�_ `RA�VC_GRP 19CdW�Q X�O�o �O�o�o�o�o�o& J1nUg�� �����"�	�F� X�?�|�c�������֏�������0�bRO�Up`I�HQP�����R��8�?T쀟3�|�����>��  Dڟl�l��@@�B�������o�4�g`SMT
mcJtm蕗�������AHOSTC]R19KO�pP�a�k M������0�  27.0zG�10�  e'� t���������b�ۿ�����4�˿ų	anonymous8� f�xϊϜϨ����л���%�'��[�0�B� T�f�x�ǿ�߮����� �Ϗ�E��,�>�P�b� ��������������� ��(�:���^�p��� �����������  $s�������� �����K� 2 DVh������� ��5GYkm7/ �v/�/�/�/�/�/ �/??*?M/��r? �?�?�?�	//-/O A?c/8OJO\OnO�O�/ �O�O�O�O�OOM?_? 4_F_X_j_�?_�?�? �__%O�_oo0oBo �Ofoxo�o�o�o�__ !_�o,>�_�_ �_��o��_��� �So(�:�L�^�p�� ��o��ʏ܏� �u�~١ENT 1LO�� P!��E�  A�3�p�_���W� ��{�ܟ���ß�6� ��Z��~�A���e�Ư �������� ��D�� h�+�=���a�¿��� ��
�Ϳ�@�/�d�'� ��KϬ�oϸϓ���� ��*���N��r�5ߖ� Y�k��ߏ��߳����QUICC0!����p�3�1q�M�_���3�2�����!ROUTER������`�!PCJ�OGa�<�!1�92.168.0�.10:��NAM�E !"�!R�OBOT���S_�CFG 1K"�� �Au�to-start{ed`tFTPkH���s��� ���$�'9 \J������ Jv!3E/Y{1/ b/t/�/�/g�/�/�/ �/?'/�/:?L?^?p? �?�?Qcu�?? O O/$O6OHOZO)?~O�O �O�O�O�?kO�O_ _ 2_D_V_�?�?�?�_�O �_O�_�_
oo�O�_ Rodovo�o�_�o?o�o �o�og_y_�_1 �o��_����� �o�&�8�J�mn�� ������ȏڏ);M _a�F��j�|����� ����֟����/�ɟ ßT�f�x�������� �!�#��W�,�>�P� b�t�C�������ο� ����(�:�L�^ϭ� ��ѯ������� � �$�6��Z�l�~ߐ� ����G�������� ����T_ERR �M��.�>�PDUS_IZ   �^����U�>n�WRD� ?��� � guest\��������������SCDMNGR�P 2NX����p��\��KM� 	P01�.14 8�� �  y��}�B�    ;����� ���߇�����������������~��\��������|���  �i  �  
����ҕ�����+��������
����l��.؋�"��luop �
dy�������&�_�GROU8�OM�� �	0�p�07��	QUPD  d��U��!TY��M�@�TTP_AUTH 1PM�� <!iPeOndan�������!KARE�L:*���K�C����VI�SION SET� ://���Q/?/ i/��/{/�/�/�/�/��/"?�/>YCTRL QM�P�v5���
��FFF9�E3.?��FRS�:DEFAULT��<FANUC� Web Server�:
Y��� A<OO*O<ONO`O<��WR_CONFI�G R<� ��?>�IDL_CP�U_PC�0��B�ȩ��@�BH�EM�IN�L���DGNR_IOG�|��S�@�NPT_SIM_�DOV[TPM�ODNTOLV >3]_PRTY)X�B��DOLNK 1SM����_�_�_�_�_��_o|RMASTE�P&|R_O_CFG"o4iUODEo6bCYCLEdo4d�0_ASG 1T<���
 o�o�o�o �o!3EWi{����k�bNUM�{�Q��08`IPC�H�o58`RTRY�_CN�0
RQ�6bSGCRN>{�Q�U�1 6ba`?bUM���p����$J23_�DSP_EN� �M�ᆀOBPROqC��LUMiJOG��1V�@Q�8G�?��{?Ń�POSRE��VKANJI_`d�
_HH��V�W�L}6h�<1�C�CL_L�@�r��H�EYLOGG+INB`���Q�P�LANGUAGE� �6�B�4 ,�>�LGW�Xf?��+����x% ���?���@���'0���`$�>MC:\�RSCH\00\��?�N_DISP YM�Ĩ�|�z��<�LOCGR�BDz��DA�OGBOOK Z�kR�P�T�X��B�T� f�x�����������v6	�<��⸥����_BUFF K1[�]� I�2�� H�S�h�d�n��ϒϿ� ����������+�"�4� a�X�j�|ߎ߻߲�����ߔ�ˀDCS }]� =��;� ��C��5Y�k�}����IO 1^�k t��� ������� ��� �2�D�X�h�z� ��������������
�0@Rdx��E^PTM  GdR2 ����0B Tfx����� ��//,/>/)Ĩ �SEV:����TYP���/�/�/ �-�RS�0��*�2��FL 1_��@��9�9?K?]?o?�?�?L�?�/TPѐ��"}ݭNGNAM���p�tU�UPS��G�I���E�A_L�OAD��G %V��%	=AR�01�?��JMAXUALRM�w��x{@AdQ:��<��C��y@C��`���Oj�lM�@̀Ҁa��k �X�	�!�p+e���OΤ,R X_C_U_�_7�|_�_�_ �_�_�_oo;o&o_o qoTo�o�o�o�o�o�o �o�o7I,mX �t������ !��E�0�i�L�^��� ��Ï�����܏�� A�$�6�w�b������� џ����������O� :�s�^�������ͯ�� �ԯ�'��K�6�o����d�����ɿ�GD_LDXDISA�0����MEMO_A�P�0E ?a+
 � ѹ%�7�I��[�m�ϑϣ�y@IS�C 1ba+ � ����'T,���
ߺ�C� .�g�Nߋߝ�߬߀� ����	���?���N� "��������b� �����;�&�_�F��� �����x����� ��7��F�| ���Z���3 W>{��p����/��_MS�TR ca-%S_CD 1d͠� m/��/|/�/�/�/�/ �/?�/3??W?B?{? f?�?�?�?�?�?�?�? OOAO,O>OwObO�O �O�O�O�O�O�O__ =_(_a_L_�_p_�_�_ �_�_�_o�_'ooKo 6o[o�olo�o�o�o�o �o�o�oG2k V�z����� ��1��U�@�y�/�MKCFG e�--��<"LTAR�M_��f��� v�����㰟METPU�n����5)NDSP_CMNT�����#�N&  g-.a�v��y���#�POSC�F/�:�PRPM�.� �PSTOL �1h��4@��<#�
��t������� ��/�q�S�e����� ��ݯ��ѯ����I��+�=��i�#�SIN�G_CHK  ~ǟ$MODAQӃ�i��a�����DEV� 	K*	MC}:�HSIZE��--ȹ�TASK �%K*%$123456789 V��hŷ�TRIG 1�jK+ lK%%�a���  ������M#F8�YP#���5$���EM_INF 1�kڇ �`)AT&FVg0E0��a�)I��E0V1&A3&�B1&D2&S0�&C1S0=P�)�ATZaߵߜ�H@����p���	��A�@9���]�D��� G� ��k�}ߏߡ����6� m�Z�l���K����� ������� ������ hs�-�����}�� ��@Rv );M_���+ /*/�N/	/r/�/k/ �/[m�/���&? 8?�\?�/�?;?E/�? q?�?�?�?O�/4O�/ �/??�OA?�O�O�? �O�?_�O_B_)_f_~��ONITORJ��G ?��   	EXEC1p���R2�X3�X4�X5��Xy��V7�X8�X9p��R0Bd�Rd�R d�Rd�Rd�Rd�R�d�Rdbdbc2�h2'h23h2?h2�Kh2Wh2ch2oh2�{h2�h3h3'h3��R��R_GRP_�SV 1��>ї�(�q�� �>Ee�S�<G���X������>c.w�@�_DR&Λ��PL_NAME �!��p�!�Default �Personal�ity (fro�m FD) ��R�R2-q 1m)d?eX)dh��q7�X dv� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V�h�t�2�������Ο������(�:���< ��d�v���������Я@�����*��R,rg 1r�yհ\��O, �����f�� @D�  z�?����f�?������A�'�6z�ܿ��;��	l��	 �xJ԰������˰ �<� ��� ���IpK�K ���K=*�J����J���JV�尻�"�ɱT���:�L�Ip@j�@wT;fb��f�n����%�4��=�N�����I��g��a�����*���*  ´  ���P�>��������n�?z��{�n���Jm���� 
�ғ�%���ت�9��� �`��  P}pQ}p�>}p|  �r�/����+�	'� �� ��I� ��  ��J�:��È��È=������6Ç�	�ВI�  �n @@
�+�l�$��l����9�A�7�N�p|�  �'��_���@2���@���f£�@֧�C��C�pC�W@ C��C��C��=o�
�A�q� "  @�U��
0�B�p"*�A��2���`�o�R�n�Dz��q��߁�������2��( �� -�����������o� ����!�o�M� �??�ff ��/|A�� ��v��7�a��
>��  P��2�(o��e������ڳڴD�?˙�o�x"Ip<
�6b<߈;����<�ê<�? <�&�K�NA둳��nO�?offf?�?&��3�@�.��J<?�`�M�� ���.ɂ�����l ƴa2//V/A/z/e/ �/�/�/�/�/�/8�F�p�/4?�/X?��y?�K?�?��E��� E��G+� F���?�?�?O'O`OKO6OoO.�BL��B�_0���OUO[� �OcO_o?5_�?\_�O��_�_�_�_U
�h�y�V�W>�r_�on_/oo,oeo�GA��d;���CRo�oNoD������o�o%�5yķD��8C|�spCH5"Z�d����a�q@I��~N'�3A�A��AR1AO�^?�$�?��;���±
=ç>�����3�W
�=�#���{e���n�@�����{�����<���~(�B�u���=B0��?����	���H�F�G����G��H�U`�E���C�+����I#�I���HD�F���E��RC�j�=z�
I���@H�!H�(� E<YD0 9ڏ�׏���4�� X�C�|�g�y�����֟ ������	�B�T�?� x�c����������ϯ ���>�)�b�M��� q��������˿�� (��L�7�Iς�mϦ� ���ϵ������$�� H�3�l�Wߐ�{ߴߟ� ���������2��V� A�z��w�������������R��q(��q�����<���e��v����a3�8������a�4Mgs������I�B+���a���{�&&	fT��x���eP�P��A�O	\���*<��R^p������  �� ��*//N/</r/��)�O� ��/�/�% �Q�/�/�/??'?9?  N?l/�?�?�?��?�?�2 F��$�Gb���A���@a�`rqC��C@��oTO�dq�|KF�� Dz@�� F?�P D��eO�O�I�cO�O�O__�1_�c?���@@*8Z^4� � �u� �n
 8_ �_�_�_�_�_�_oo +o=oOoaoso�o�zuQ� �����1���$MSKCFM�AP  R5� `6uQqQ��n�cONREL  ��a� �bEXCFENBwq
�c�e qFNC'�tJOGOVLI�Mwdprd�bK�EYwsu�bR�UNc|su�bS?FSPDTY�p)v<u�cSIGNt�T1MOTeq��b_CE_GRP� 1sR5�c\ :�I�2�m���Di��� a�Ώ��Ï���(�ߏ �^������K���o� ܟ��ɟ�H��� l�~�e���Y�Ưد������F�`TCOM_�CFG 1t�mЀV8�J�\�
�_A�RC_$r�2yU?AP_CPL��6t�NOCHECK {?�k � ׸տ�����/�A� S�e�wωϛϭϿ�������kNO_WAI�T_L�w�e�NT� �u�kw[5�_7ERR!�2v�i�� ߠ߲߾���c���ߴ�T_M�Oc�wj�, ��B�3���PARAuMd�x�k�tV`#���=?�� =@�345678901������������ +�U�g�C�����y�觃�����t���U�M_RSPACE��olV>H�$OD�RDSP��v2xO�FFSET_CAsRT��yDIS��yPEN_FIL�E� jq^�+�v�OPTION_IO��YPWORK 5y'�5s x��fRuQ��2��2	C �	2��[ �RG_DSBL  R5sx\�zRIENTTOp!C�oP�a.A[ �UT_SIM_D���b�b[ V_ LCT z?�*+�^�)�_PEXE�,&RAT8 jv2u��p0"� UP {.�PS0��/�/�/��/�)�$O�2 �m�)deX)dh�>�X d��? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�H2
?�O �O�O�O�O__1_C_U_%�<�O_�_�_�_ �_�_�_�_o!o3oEo�O� �Ov 1r(?���(��0}7�, �l�p�` @D�  &�a?��c�a?m�a�%�D�c�a���l;��	l�b	 �xJ�`�o�u��` ��< �	p� ��r��H(��H�3k7HSM5G��22G���G�p
�������XYk|��CR�>�qȋs�a����*7  ���4�p�p���pT���B_����j%���t�q� �)�/��aD������_6  ���P� UQ� �� |Б��������	'� �� ͂I� ��  ��i�=��������a	����I  �n @)��mC���"m��[��N����  '� ��~q�pCN�C�@�s�pC�t��ҟ 5�
��*=x@#�7~9�^�n�B�I�A��Q���G 0�q��bz毀�������ȯ�����( �� -݂*�΁6���AFm� �0rx��m�~lp �?�ffU ܫN�`�����n�8m྿̺>�  P�aզ(m�������� q�c�d#?˙�m�xA�n�<
�6b<߈;����<�ê<�? <�&1jςm�A0��c���n�?offf?0�?&�����@�.�J<?�`��l�� ���dѩ�e�ϟgߋ� �d��Q�<�u�`ߙ߄� �ߨ��������)� � M�8�q���
��j���~f�E�� E�0�?G+� F���� ��� �F�1�j�U���(y�[bB��A��|� ���t�z���3�� T��{�������t��h��u�w�>��*�N9K���A��Z�_��Cq�mc��?Ƀ�//D///T)����pٞ�a�`CH�T/A
$� !�!@�Iܝ�'�3A��A�AR1A�O�^?�$�?������±
=�ç>����3�W
=�#�>���+e�� �������{����<���.(�B��u��=B0�������	�3�\*H�F�G����G��H��U`E���C��+�Y-I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0X/�?O�?/OO SO>OwObO�O�O�O�O �O�O�O__=_(_a_ s_^_�_�_�_�_�_�_ o�_ o9o$o]oHo�o lo�o�o�o�o�o�o�o #G2kVh� �������1� C�.�g�R���v����� ӏ��Џ	��-��Q� <�u�`�������ϟ�� �ޟ��;�&�8�q�:\�(����,������]���x����p!3�8���<ӯp!4Mgs�����IB+�+��a?���{�E�E����s�����Ϳ���Pe�P��(�{�`4��I�[�իR}�����ϳ�������  ���˿I�7�m�[� ���H� ߿�����������"�4�F�X�  m�ߵ����������2 wF�$�Gb���²����!C����@�s����� F�� Dz/��� F�P D�����������,>P�?��ͫ@@W
}���ԉ������
 W���� &8J\n�����*� ���˨��1��$PARA�M_MENU ?�q�� � DEF�PULSE�	�WAITTMOU�T+RCV/ �SHELL_�WRK.$CUR�_STYL �G,OPT]�]/PT�Br/l"CB/R_DECSN ��,�/ �/�/
???)?R?M? _?q?�?�?�?�?�?��USE_PROG %�%�?#O�3CCR ��6G�_HOST !F�!;DxO0JT�BO�C[OmA�C�O/K_TIME"�B��  �GDEB�UG�@��3GINP_FLMSK�O�(YT��9_*UPGA�UP \��g[CH�6_'XTYPE����?�?�_oo#o 5o^oYoko}o�o�o�o �o�o�o�o61C U~y����� ��	��-�V�Q�c��u���*UWORD �?	{]	RS���	PNSW��V$ڂJO�!��T�E�@�VTRACE�CTL 1|q��� �� ���4��_DT Q}q�c��(�D � � y� �Rp�-t�p�.��/��U0��1��2��3��U4��5��6��7��U8��9��:��;��U<��=��>��?�� n ��]���� ��� ��D��Z ��F��P��H��I��J���P��EL��M��� ��O�����Q������ဆ�T ��U��V��W��UX��Y��Z��[��U\��]��^��_��U`��a��b��c��Ud��e��f��g��Uh��i��j��k��Ul��m��n��o��Up��q��r��s��Ut��u��v��w��x��s����� ��� ����P��� ��� �������	��
���������������@�������������V���*����������(��� ������ਆ�N���!��"��#���'���%��&��'���(��)��*��+��,����������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿոl�x��� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_x� ���_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� ��_@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/�L/^/h!�$PGT�RACELEN � g!  ���f �|&_�UP ~��e��!� �!� �|!_CFG ��%�#f!� ���$� �/�/;�"DEFSPD ��,�1�� �| IN~� TRL ��-�f 8�%G1PE__CONFI� ��%���!�$�<LID�#��-~�4GRP 1��7�!�g!A ����&fff!A+�33D�� D]�� CÀ A@6B1�f d�$I&I��1�0� 	 p?�"�+@O ´yC[ODKB|@�A�OmOO�O�O�Of!>�T?�
5�O4_F^0_� =��=#�
K_�_G_�_�_�_�_ �_c_�_&o�_6o\oGo�  Dz�c�of 
 qo�oao�o�o�o�o 0T?xcu������IK
V�7.10beta�1�$  A��E/�ӻ�Ay f ,�?!G�C�/>��+���0T����+�BQ�c�A\i�T�D;�{�p�"�B������Ə؏�T�O'O�2�8��\�G���k� ������ڟş���"� �F�1�V�|�g����� į���ӯ���	�B� -�f��ov���K����� �������>�)�b� M�rϘσϼϧ�����<�=�F@ �� '�۫%Wك�W߉ߛ� �6���������%� �I�4�m�X��|�� ����������3�� W�B�{���x������� ������S~� w�8����� �+O:s^ ������
�<�/ /R�d�v�l/~/�ߥ/ ��������/�#?5?  ?Y?D?}?h?�?�?�? �?�?�?�?O
OCO.O gORO�O�O�O�O�O�O �O	_�O-_?_jc_u_ $_�_�_�_�_�_�_�_ oo;o&o_oJo�ono �o�o��(/�ob/ P/&Xj�/��/�/ �/�/��o��3�E� 0�i�T���x�����Տ ��ҏ���/��S�>� w�b�������џ���� ���+�V_O�a���� p�����ͯ���ܯ� '��K�6�o�Z����o �o�o޿*<n D�rk�}Ϩ��� �φ������
�C�U� @�y�dߝ߈��߬��� ������?�*�c�N� ��r��������� 0���;���_�q�\��� �������������� 7"[F����ο ����(�0^� Wi�Ϧϸ�v�r ��/�///S/e/ P/�/t/�/�/�/�/�/ �/�/+??O?:?s?^? �?�?�?�?�?�?�O 'O�?KO6OoO�OlO�O �O�O�O�O�O_�O_ G_2_k_����_�_ �
ooJCoUo ����oL_�o�o�o �o�o?*cu `������� ��;�&�_�J���n� ����ˏݏO�� 7�"�[�F����|��� ��ٟğ���!��� W��_�_�_�����_�_� o���6b�$PL�ID_KNOW_�M  bd��j�#�SV ��3e=�:e��z�����7��¿������j�vmC�M_GRP 1�P���`d�bd@I�߶B�_�
�_��� ��t��@ǘϾ�^��� �ϮϪ�
�����F�� d�(�Zߠ�^����ߔ� �����*��� �f�$� L��Z�|���������,�>�#�MR'Éb.�Tg��� � ���������������� ����Q+%7�� �������� M'!3��������Y�ST'�1W 1�3e3 �i�;0:o A >/g� </N/`/r/�/�/�/�/ �/�/�/?C?&?8?y? \?n?�?�?�?�?�?	O�'2(.:/j��	<=O.3'O9OKO]O�!#4vO�O�O�O!#5 �O�O�O�O!#6_&_8_J_!#7c_u_�_�_�!#8�_�_�_�_!#M_AD  wd3#�x`$PARNUM  ++�5o"WSCHOj ]e
�gppa�i=��eUPDpo��e�t"_CM�P_$�R`ؠ`'�;�)tER_CHK7u��;�Or4F{�RS|�2�#�_MO�Q`��u_�be_R/ES_G' �+-O ���H�;�l�_��� ����Ə���ݏ����w&@�|�5��u u@R�q�v��s�@���� ���sPП����sbP �.�3��s�PN�m�r���s `�������rV �1�P���b@cX���p�$@cW��(��(�@@cV��4���rTHR_�INR|�Taud�<�MASSI� Z�]�MNH�{�MON�_QUEUE Q�.�bvg��g�bdN.pUrqN��`{ΰ�ENDб��EX1E����`BE��ڿ>˳OPTIO׷�{�ΰPROGRAM7 %��%Ͱ���o̲TASK_I�Qd@�OCFG Ꭾ��o����DATuAe���@�2�N�`�r߄ߒ�<� �������ߖ��!�3�xE�W�
�INFOe��"ݘ������� ������)�;�M�_� q����������������n�z�"� �!���OpDIT ���s�WERF�L��#RGADoJ �b
A��0��?��P��IOORITY��av��MPDSPX��eU����OG$ �_TG� K���ET�OE��1�b _(!AFD�E�p���!tcp|��!ud�>�?!icm��nFXY_���b{���)� *J/\/` ���G/�/k% w/�/�/�/�/�/?�/ 2??V?h?O?�?s?�?z�?*�PORT3��Rc���u�_CARTREP�|bk@SKSTA��^�zSSAV���b
�	2500H8�63(�ς5D1�*b`@�����s�O�O�G	PURGE��B�	�yWF�@DO��$�evW�T�a��:WRUP_DE?LAY �bT�R_HOT{��%�o�_TR_NOR�MAL{�}_�_�VS�EMI�_�_oCaQ�SKIP1��u�Cx 	bO\o\@ Jo�o�o�ojh�u�o�g �o�o	�o?-O u��_���� ���;�)�_�q��� I�������ݏ��Ǐ %��I�[�m�3�}������ǟٟ�ͥ�$R�BTIFR�RCgVTM.+D�	��DCR1c�8l����C���D�OC�T�?�(�p?9!w<!\�!em�&�$�F���¼詿��߿����eo���o <�
6b<߈;�܍�>u.�?!<�&ǯ ���)�ŰHB�T�f� x���������ҿ��� ���>�)�b�Mφ� qσϼϟ�����5�� (�:�L�^�p߂ߔߦ� �������������6� !�Z�E�~��s���� 	������ �2�D�V� h�z������������� ��
��.RdG ������� *<N`r�o �����/�&/ 	//\/��/�/�/�/ �/�/�/�/?"?4?F? X?C/|?g?�?�?�?�? �?�?�?O0Os/TOfO xO�O�O�O�O�O�O�O __,_OP_;_t___ �_�_�_�_�_�_oGO (o:oLo^opo�o�o�o �o�o�o�o�_�_$ H3lW���� �o�� �2�D�V� h�z�������ΈB��GN_ATC 1��O� AT&FV0E0΋�ATDP/6�/9/2/9��ATAΎ,�AT%G1%B9�60�+++�3�,.�Hc�,B�I�O_TYPE  �����ЏRE�FPOS1 1�>�� x��������?�P���� 6�������V�߯z��� �9�Ǜ2 1�����$��� �ƿ<D�ё3 1�^�p������:�%�^�ܿS4 1����Q��������q�S5 1� �ϚϬ���d�O߈��S6 1��/�A��{�������S7 1���������y�|��0�S8 1�G�Y�k��#��G���SMASK 1����  
����e�XN	O��;�A�����͑?MOTE  ��ʔ���_CFG ������̒PL_RA�NG���q��POW_ER ��^ ���SM_DRYP_RG %��%����dTART ��V�
UME_P�ROs� ʔ_E�XEC_ENB � =���GSPD�� #��4TDB�>PRM_PMT�_m�TQ ����O�BOT_NAME� ���׉O�B_ORD_NU�M ?V���H863  ��t ���!\<�  # w	r*!@�"�D|<���PC_T�IMEOUT6 �x��S232
1��� LT�EACH PEN�DAN_ ����e����Main�tenance �Cons�r���*"��/�KCL/C�� :���/? �No Use�e��/U?�v#NPO�218�����t!CH_L� ����7�	�1�;MA�VAIL�a#����t!PACE1 ;2�ٜ �?% dH�9�eF%�<�>�L8�?H �9 �O�?�O�O_�O(_#W TOfOxO�O8_�O�O�_ �_�__o i��4m T_f_x_�_�_�_�_�o �o�oo .�5;A2@NROdovo�o6 �o�o����4��I�N{3]o��� S������ޏ0�Q�8�f�N{4z������� p����8���M�n�U���N{5������ ͟ߟ���%�4�U�� j���r���N{6��Ư د����� �B�Q�r�@5χϨϏϽ�N{7ѿ �������=�_�n߀��Rߤ��߬���N{8 �� ��$�6���Z�|� ���o���������N{�G ��� t���$
�� C� e#p������������� :hL���2��+��^�!dt Y�k���� �����8o R~q���� ��//=/7I km�/���/�/�/ ??+?=?3/]?W/i/܋/�= `�� @NP�5<�?�/�) A�5�?1OCOI?#J$O VO�O�O�O~O�O�O_ �O�O�O_^_ _2_D_ v_�_�_�_�_�_o$o��_�_
o<o~o@oN<
�O�oN{_MODE�  +��iS E�+��ox?v:_��?'y�z	��o��CWORK_AD��m��q�R  +�����p_INTVAL�`�@�zR_OPT�ION1� u���VAT_GRPw 2�+�]�G(���L�� ԏ揥�
��.�@� ��d�v���O�o���d X�ß����ϟ1�C� U�g�)���������ӯ �{�	��-���c� u���I�����Ͽ�� ϛ��;�M�_�!σ� �ϧϹ�{������� %�7���[�m��Aߏ� �����ߛ����!�3� E�W���{����s� ���������/�A�S� e�w������������ ��+��Oas ���?��� �'9K[�����e�$SCAN�_TIM�a��\���R �(�3�0(�L8z�W�p�p
Wt�Z��2#Nq!�#�Y�:.(/1�#"M"2{$!!d�(~!"�!�r #])�0���/�/�/�r�)�/  �P5�0�2 � 8�?U?g?>1D��j?�?�?�?�? �?�?�?O#O5OGO?Nq�%RO�O�O�[N![q;�o�t�Nqp]M�t��Di�t!c{  � lM"Nq�A !
%�1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�gS�o�o�o '9K]o��� ������#�5� G�Y��o�o�K������ Џ����*�<�N� `�r���������̟ޟ�����1�  0 �B|�_g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ �p���)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� ���ϐ�������� �0�B�T�f�x��� ������������,�0>�P�J�V�  �1�� �������������� 1CUgy��������	 �y3"HZl~ �������C&a5/</+&�r!� 5/q-	12345678R_���L{0�@�/�/�/�/�/?3,?>?P?b?t?�? �?�?�?�?�?'OO (O:OLO^OpO�O�O�O �O�O�?�O __$_6_ H_Z_l_~_�_�_�_�O �_�_�_o o2oDoVo hozo�o�_�o�o�o�o �o
.@Rdv �o������� �*�<�N�`������ ����̏ޏ����&� 8�g�\�n����������ȟڟ����"�+& s�C�U�:�Z���������Cz  Bp�   ���2�/$@��$SCR_�GRP 1�(��e@(�l��� @ >Z! U!m��	  #�-�=�6�n�p�l�S��y(J�w�e������3%Dʰ֠o���ป��M-�10iA 890ƅ%90� Ɓ M61C �#�-I���*#�
\�l�,�O'�|�Z!�S�;�o�}�	�n�����������X �,���Y"N�a� ���ߖ�i�@�.!`/���m�����"��B�BŠ�J�H�a�H�A֠p�  @. ��l��?���D�HŠ����H�F@ F�` �������;�&�K� q�\�������<���`��������B� ��YD}h��� ����
CҾ�?4#��0/v/�%��
��������V��j�@���/ B�*'��P����EL_DEFAU�LT  C�����X!M�IPOWERFL�  P�p%W"} W7FDOe& p%���ERVENT 1O���I�n#=��L!DUM_E�IP��(�j!?AF_INEd ?��!FT�/7>��/[?!K߀? ��J?�?!RPC_OMAIN�?�8��?��?�3VIS�?�9���??O!TP2@P�U6O�)d.O�O!
�PMON_PROXY�O�&ezO�ORB�O�-f�O#_!R�DM_SR��*g_o_!RL(�_�$Yh^_�_!
�0M�O��,i�_o!RL�SYNCo.i8|�_So!ROS�/zl�4Bo�on?�o2S �o�o�o�o5�oY  }D�hz�� ���1�C�
�g�.����R����'ICE_�KL ?%�+ �(%SVCPRG1��������3$�)��4L�Q��5t�y��6����뀁7ğɟ�=��/�9��脆_A��� i������>���� f��끎�	�끶�1� �ޟY������.� ���W�ѿ����� ��!��ϯI����q� �����G����o� ���������9�;� 翹�˂�ҏ䀄��� á������� �9�$� ]�H���~����� ������#��5�Y�D� }�h������������� ��
C.gR� v�����	� -QcN�r� �����/)//�M/��_DEV ��)�MC:�U(��]g$OU�TYB`!x&c(RE�C 1���` � � `  	 *` ` ` ` �!��!U+�#��U/�.D�$`!�"?`!)A�8�+
 �P�b�6 s�'�  �  '� ��    Cf���"�#�!� U` /` �` ��=�y �y �y ���+��` B� D�?O�%��|0��<S  M��H� �0_�k�? O�` ��4)` ��?��T`!y ��0�` k� �NPO�OOc݀;�[0�0�1o  k�=0i�O !� U� �` ` ,` -�xO��y ��!�D�n� M�O]_�Oc��O�@�F��O
__�._@_R_d_If�6r _�H�i@_0�2��x�C�@��_�!er` �\4�P#�_��fy �y �y ��y �` To�ooh}$0k �  � ~�1   �i@�=�o ;@�2�0 l` K`$|o�dy %�y �y Dq��! ,a�oh[�l�0k`��bR  Ȣ l�P
5�2` �` �V(�c�4��D��!ج�ta��; L�  "Ɣ3G�Qݢ �>` �`�� e&` ` w�F���b�D֔DX� >XX��� �aĀ<Đ?g���?�?�?�?���ď"F �;  K#f�4���'�W��  =� �� ��
j` Q� ,���y U�y �H��` U|�b�t��"x1 � �T� B�x�f�������ү�� ����,��P�>�t� ��h�����ο��޿� �(�
�8�^�Lς�p� �ϔ����Ͼ� ���$� �4�Z�H�~�`�rߴ� ���������� �2�� V�D�f�h�z����� ����
���.��R�@� b���j����������� ��*<`N��r�����%V �1��, P 8g@.�[1#�'�p^� �p(a*TYPE��/e"HELL_CCFG���&� �66�0-RS�p�� �//?/*/c/N/�/ r/�/�/�/�/�/?�/�)?8;�p:>����` %K?y?�?F=J1J1`�p�>�1�p���a22!�d�?�?�H/K 1���a�? AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_|OMM� ���_FTOV_ENO�n�wOW_REG_�UI�__IMWA�IT�Rq�6kOU�Tf iTIMne��ZoVAC�|1o#a_UNIT�S��fwMON_AL�IAS ?e�Y ( he�o�o 0��o]o� �>������ #�5�G�Y�k������ ��ŏ׏������1� ܏B�g�y�����H��� ӟ���	���-�?�Q� c�u� �������ϯ� ����)�;��_�q� ������R�˿ݿ�� Ͼ�7�I�[�m��*� �ϵ����τ����!� 3�E���i�{ߍߟ߱� \�����������A� S�e�w��4����� �����+�=�O��� s���������f����� '��K]o� ,������ #5GY}�� ��p��//1/ �U/g/y/�/6/�/�/ �/�/�/�/?-???Q? c??�?�?�?�?�?z? �?OO)O�?:O_OqO �O�O@O�O�O�O�O_ �O%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3o�_Woio{o�o�oJo��o�o�o�o�c�$�SMON_DEF�PRO ����4q �*SYSTE�M* . "vR�ECALL ?}�4y ( �}!�xyzrate �61=>desk�top-b25t�4o0:10168 ��q�q����y}
tw ���4�F�X��us�5916�'���ʏ܏o�1}�����2�D�V��w�7copy md�:program�_1.tp vi�rt:\temp\���,���ϟ�t� ����;�M�_��� ��(���˯ݯ😯�� ��7�I�[�n�����$�е�ǿٿ�t;t�fr�s:orderf�il.dat��mpback���/��A�S��z2t�b:*.*	���'ϸ���l���q6x��:\}π�������<�N���7��a����,߽��� b�t����ߪ�;�M�_� �ύϨϹ�����p� ����7�I�[��ρ� ��$ߵ�����l�}��� "�3EW�|��  ���h����/ AS�x
.� �������=/O/ b���/*/�/�/�/ r���(�9?K?]?�� ??&��?�?�?n� ��5OGOYO���?O �/�O�O�Oj/|�/�O 1_C_U_��/_�_ �_�_�Ox/
_�_�_?o Qo�_�Oo�o,o�o�o b_t_�_�o�o;M_ �_�(���po ���7�I�[��o  $���Ǐُl��� ��3�E�W���� � ��ß՟h�������/� A�S��/�/�?�.��� ѯd?v?���?��=�O��`��$SNPX_�ASG 1�������� P 0 '�%R[1]@1�.1`���?�j�% ��ֿ����ݿ�0�� :�f�Iϊ�m���ϣ� ����������P�3� Z߆�iߪߍߟ����� �����:��/�p�S� z������� ��� 
�6��Z�=�O���s� ������������  *V9z]o�� ���
��@# JvY�}��� �/�*///`/C/ j/�/y/�/�/�/�/�/ �/&?	?J?-???�?c? �?�?�?�?�?�?O�? OFO)OjOMO_O�O�O �O�O�O�O�O�O0__ :_f_I_�_m__�_�_ �_�_�_o�_oPo3o Zo�oio�o�o�o�o�o �o�o:/pS z����� �� 
�6��Z�=�O���s� ��Ə���͏ߏ �� *�V�9�z�]�o����� ���ɟ
����@�#��J�v�Y�r�PARAoM ����_ �	�z�P���j�OFT_�KB_CFG  �����ѤPIN_�SIM  ��Ʀ�)�;�ɠr�RV�QSTP_DSB� �Ƣw�����SR� ��� & �������ΦTO�P_ON_ERR�  ����P_TN ���AݲRIN�G_PRM� ���VDT_GRP� 1����  	ʧ��\�nπϒϤ� ����������%�"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�w�t� �������������� =:L^p�� ���� $ 6HZl~��� ����/ /2/D/ V/h/�/�/�/�/�/�/ �/�/
??.?U?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o Fomojo|o�o�o�o�o��o�o�o30ѣV�PRG_COUN�T����^rENB)�YuM�s㤐_UPD 1��8  
G��� ��'�"�4�F�o�j� |�������ď֏���� ��G�B�T�f����� ����ןҟ����� ,�>�g�b�t������� ��ί�����?�:� L�^���������Ͽʿ ܿ���$�6�_�Z� l�~ϧϢϴ��������VuYSDEBUG�hp�p���d�y�S�P_PASShu�B?.�LOG ���u�s������  ��q��
MC:\Z�
�[�_MPC`��u���ߒ�q��� �q��S_AV �c���l������SV��TEM_TIMEw 1��{ (�pպ�t�����T1?SVGUNS�piu�'�u���ASK_OPTIONhp��u�q�q��BCC�FG ��{I� qB��5�`5� ;zC�l�W�i������� ��������2D/ hS�w���� �
�.R=va������� �/��B/-/f/Q/ �/�/�� �/�/�/ �/�/ ??D?2?T?V? h?�?�?�?�?�?�?
O �?O@O.OdORO�OvO �O�O�O�O�O_�H� _,_J_\_n_�O�_�_ �_�_�_�_�_o�_4o "oXoFo|ojo�o�o�o �o�o�o�oB0 Rxf����� ����>�,�b�_ z�������ΏL���� �(��L�^�p�>��� ������ܟʟ�� � 6�$�Z�H�~�l����� ��دƯ��� ��D� 2�T�V�h�����¿x� ڿ�
��.Ϭ�R�@� bψ�vϬϾ��Ϟ��� ����<�*�L�N�`� �߄ߺߨ�������� �8�&�\�J��n�� ����������"�ؿ :�L�j�|�������� ������0��T Bxf����� ��>,bP r������/ �//(/^/L/�/8� �/�/�/�/�/l/? ? "?H?6?l?~?�?^?�? �?�?�?�?�?OO O VODOzOhO�O�O�O�O �O�O�O_
_@_._d_ R_t_v_�_�_�_�_�/ �_o*o<oNo�_ro`o �o�o�o�o�o�o�o 8&\Jln� ������"�� 2�X�F�|�j�����ď ��ԏ֏���B��_ Z�l�������,�ҟ�������,��J��$�TBCSG_GR�P 2����  �J� 
 ?�  u� ��q�����ϯ��˯���)�;�N�U��\�_d, �j�?J��	 HC��8�>�����9�CL � B�m�����z���β\)��Y�  A���B��;��Bl�=�,�����Z�,��  D	 �{�F�`�j�Cs���H�Ϧϰ̖���@J� �+�>�Q��.�|ߙ�@d�v��������؈J��	V3.00~m�	m61c��	*,�$�I�;�D�>���J�(��� qr�D�s�  #�����D���N�J�CFG ��ef� i������������� �7�E��E�k�V��� z��������������� 1U@yd�� �����? *cN`���� ��m����/"/� U/@/e/�/v/�/�/�/ �/�/	??-?�/Q?<? u?`?�?�?J�6��?� �?�?�?*OONO<OrO `O�O�O�O�O�O�O�O __8_&_H_J_\_�_ �_�_�_�_�_�_�_o 4o"oXoFo|o�o���o �obo�o�o�oB 0fTv���~ �����>�P�b� t�.���������̏Ώ ����:�(�^�L��� p�������ܟʟ �� $��4�6�H�~�l��� ��Ư���د�� ��o 8�J�\����z����� ���Կ
���.�@�R� d�"ψ�vϬϚϼ��� ������<�*�`�N� ��rߨߖ߸ߺ���� ��&��J�8�n�\�~� �������������  �"�4�j�X���|��� ��n���������0 TBxf���� ���,P> t���d��� �/(//L/:/p/^/ �/�/�/�/�/�/�/?  ?6?$?Z?H?j?�?~? �?�?�?�?�?�?OO  OVO��nO�O�O<O�O �O�O�O�O_
_@_._ d_v_�_�_X_�_�_�_ �_�_o*o<o�_oro `o�o�o�o�o�o�o�o 8&\J�n �������"� �F�4�V�|�j����� ď������O�$��O ��f�T���x������� �ҟ��,����b� P���t�����ί௚� ����(�^�L��� p�����ʿ��ڿ �� $��H�6�l�Z�|�~� ���ϴ��������2�  �B�h�Vߌ��8��� ��rߠ�����.��R� @�v�d������� �������N�`�r� ��>�������������  J8n\� ������� 4"XFhj|� �����/0/�� H/Z/l//�/�/�/�/ �/�/�/??>?P?b? t?2?�?�?�?�?�?�>�  @
C �
FO
B�$TBJ�OP_GRP 2���5�  ?�
G6B=C��DL��0�xJ�@��
D@ �<� ��@�
D �@@UB	 �C��� �Fb  C�xVGUAUA>����E��E�I>��@�A�33=�CL�@�fff?�@?�ffB�@Q�E-_8W�N���O>�nR�\)�O�@�U����;��hCY�@��  @�@UAB� � A�$_�_�S�UC�  D�A�LwP��RO�z_�Sb���
:���Bl�P��P�D�Q�_So
A?Aə�A�hcZQsDXg�F�=q�e�
o�@�p��b�Q�;�AȰ@�ٙ�@L�CD	�x`�`�o�ojo|o>BÏ\u�oh�Qts}�a@33@QV@C��@�`ew�o>��D�u*�@�� p�qP<{�Nr�@@�PZv_p�� ��&�:�$�2�`��� l�&���ʏ����!� ����@�Z�D�R������DT�
Fґ�E	�V3.00�Cm761c�D*���D�A
�� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,I&�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^'`;Q���8�E`F�O���
F���Q��K�2DES�TPARS  ��8O@3CHRe�AB_LE 1�DK.�
CP�%� ~ �P��P�P�	GAP�	�P�
P�P���
A�P�P�P�|�RDI��NA����¿Կ���`�Oh�z˄� �ϨϺ��΀�Sf�LC *ʍߟ߱������� ����/�A�S�e�w� ���������)Me� iߘ�$���1�C�￀��%�7�IȀ�
�N�UM  �5*NA�@@ ��[����_CFG ������A@6@IMEBF_TTk���LCx�5VERY�6�K�5R 1�DK
' 8�
B@� �0/�  ��� ���� 2D Vhz����� /�
/S/./@/V/d/�v/u_��b@L
�6@MI_CHAN�A L �#DBGLVPCL5A� �ETHERAD �?�550�M���/�/N?0F� ROUmT_ !DJ!�4��?q<SNMASK�*8LC;1255.��5��?�?2DOOL�OFS_DIk���%9ORQCTRL �mK���hM8WO�O�O�O�O�O�O �O
__._@_�|ON_�`_�_a�PE_DE�TAI8-JPON?_SVOFF#O�S�P_MON ��J�2�YSTRT�CHK �DN�g?�RVTCOMP�AT�X53�T�PFP�ROG %DJ%}	qaRAM_17o<�\APLAYl��Z_INST_M�0e �l�W�dUS_�WoibLCK�l�kQ?UICKME� #�ibSCRE@p>-:tps�ib �a[p`y�"qp_uy���Ti9SR_GRP� 1�DI ؕ�0��z�� �5�#�Y�G��2 �� ��S��o����܏ǅ�� ��)��M�;�q�_� ������˟���ݟ���7�%�G�m�	1?234567堃����b�XZu1��{
� �}ipnl�/ՠgen.htm�����*�<�R��Panel _setup@�}6o���������ȿڿ  o�e��$�6�H�Z�l� 㿐�ϴ��������� ߅ϗ�D�V�h�zߌ� ���C�9�����
�� .�@��d��߈��� ������Y�k��*�<� N�`�r��������� ������8��\�n����-�nU�ALRM�`G ?=DK
  � 	L?pc�� �����//6/~�SEV  ��h&�ECFGG ��]�&��A�!�   Bȣd
 7/�c-5�/�/�/? ?%?7?I?[?m??�74t!�r��[ �3ȏ��?B'Imf?wk�P(%*/O`
OCO.OgO RO�OvO�O�O�O�O�O`	_�O-_�<�d �=��?;_I_?pHIS�T 1��Y  �(�  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupage,153,�o��_�_oo �� �_�]936�_lo~o �o�o1b�o�o�o�o %�oI[m� �2�����!� �E�W�i�{������� @�Տ�����/����S�e�w���������� L��QL������1� C�F�g�y��������� P����	��-�?�ί �u���������Ͽ^� ���)�;�M�ܿq� �ϕϧϹ���Z�l�� �%�7�I�[���ߑ� �ߵ�����ğ֟�!� 3�E�W�i�lߍ��� ������v���/�A� S�e�w���������� ������+=Oa s������ �'9K]o� �������� ��5/G/Y/k/}/�/� �/�/�/�/�/?�/1? C?U?g?y?�?�?,?�? �?�?�?	OO�??OQO cOuO�O�O(O�O�O�O �O__)_�OM___q_ �_�_�_6_�_�_�_o o%o/"/[omoo�o �o�o�_�o�o�o! 3�o�oi{��� �R����/�A� �e�w���������N� `�����+�=�O�ޏ s���������͟\�����'�9�K�6o���$UI_PANE�DATA 1�������?  	�}]���`��ȯگ��� ) � $�ᔒ�O�a�s����� ���Ϳ�����'� �K�2�oρ�hϥό������������ Ha$�7�<�N�`�r� �ߖ��Ϻ�-������ �&�8�J��n�U�� y����������"� 	�F�-�j�|�c�������������� +=��a�߅�� ���F�9  ]oV�z�� ���/�5/G/�� ��}/�/�/�/�/�/*/ �/n?1?C?U?g?y? �?�/�?�?�?�?�?	O �?-OOQOcOJO�OnO �O�O�O�OT/f/_)_ ;_M___q_�O�_�_? �_�_�_oo%o�_Io 0omoofo�o�o�o�o �o�o�o!3W> {�O _�_���� ��pA��_e�w��� ������&����܏�  �=�O�6�s�Z���~� ��͟���؟�'�� �]�o���������
� ۯN����#�5�G�Y� k�ү��v�����׿� п���1�C�*�g�N� �ϝτ���4�F���	� �-�?�Qߤ�u߇��� �߽��������l�)� �M�_�F��j��� ����������7��[�����}�l�������������)��$�� Pbt��� �����(L 3p�i������ /(�����$U�I_PANELI�NK 1����  � � ��}1234567890Y/ k/}/�/�/�/�$��W/ �/�/??+?=?�/a?�s?�?�?�?�?S9S h*�=��U   �? O(O:OLO^O�?\1O �O�O�O�O�O�O�O_ (_:_L_^_p__~_�_ �_�_�_�_�_�_$o6o HoZolo~oo�o�o�o �o�o�o�o
2DV hz$�����
�E0,/A�M� /�p�S�������ʏ܏ �� ��$�6��Z�l� O����<�?�����T! ���1�C�U�g�Z3 ��������ǯٯ�z� �!�3�E�W�i��<�� ������C��ÿտ� ���Ϥs5�G�Y�k� }Ϗϡ�0��������� �߮�C�U�g�yߋ� ��,���������	�� -��Q�c�u���� :���������)��� M�_�q���������(� ����~���7I, mb����� ��3ƞ����՟ w��������/ ��,/>/P/b/t/�// �/�/�/�/�/??�� ����^?p?�?�?�?�? ?��?�? OO$O6OHO �?lO~O�O�O�O�OUO �O�O_ _2_D_�Oh_ z_�_�_�_�_�_c_�_ 
oo.o@oRo�_vo�o �o�o�o�o_o�o *<N`���� �������8� J�-�n���c�����ȏ ڏI��m"��F�X� j�|��������/֟� ����0���T�f�x� ������?/?A?�o� �,�>�P�b��o���� ����ο�o���(� :�L�^�p����Ϧϸ� ������}��$�6�H� Z�l��ϐߢߴ����� ���ߋ� �2�D�V�h� z�	����������� g�.���R�d�G��� k������������� ��<N1r�� ��;��&8 J=�n����� �i�/"/4/F/X/ ǯٯ믠/�/�/�/�/ �/?�/0?B?T?f?x? �??�?�?�?�?�?O �?,O>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_#_�_ �_�_�_ oo$o�_Ho Zolo~o�o�o��o�o g�o�o 2Vh K�o���������o�/�/�u���$UI_POST�YPE  �%?� 	e������QUICKMEN  ��d������RESTORE �1ݏ%  ���,�>�b�m]��������� Οq����(�:�ݟ ^�p�������Q���ů ׯI��$�6�H�Z��� ~�������ƿؿ{��� � �2�D��Q�c�u� 翰��������ϛ�� .�@�R�d�߈ߚ߬� ����{υ����s�%� N�`�r���9���� �������&�8�J�\� n��{���������� ��"��FXj| ��C����ނ�SCREր?�ۍu1sc�'�u2G3G4�G5G6G7G8<G��USER).2@T(IksQ�U4�5�6�7��8���NDO_C�FG ޖ�  �&� ��PDAT�E ���None V��S�EUFRAME � ��&!RTOL_ABRT1/���H#ENBR/C(G�RP 1���?Cz  A��#�!���/�/�/�/�/ 6
??A*ՀUr(A!a+?MSK  u%}1�a+N.!%[�~2%���?��VISCA�ND_MAXs5�I�](�0FAILO_IMGs0`����#}(�0IMREG�NUMs7
�;BS�IZs3&����,CONTMOU4Q u4��PE�_�c�� �@��"�FR:\�? �� MC:�\RC\LOG�FB@� !�?�O�A��O_�z �MCV�O�CUDM1*VEX3[�`�TqF�"ᖉ�`(��o=��͍_��Z �_�_�_�_�_�_�_o o,o>oPoboto�o�;_PO64_9C�B Κ�n6�eK LI�A�j�h�aV��l�f@�g�o� =	��hSZV�n�����gWAI�o�4ST�AT �+�@�O���z$���5�J!2DWP  ��P G)����a��;@'��2_JMP�ERR 1㖋
�  ��2345678901|����� ��ď��ɏ���� B�5�f�Y�k����<N0MLOW{~�@�0�@g_TIYH�'�0�MPHASE  �%���3SH�IFTO21"x[
 <���?\��;� a���q���Я����� ݯ��N�%�7���[� m�������ɿ�ٿ뿀8��!�n�E������*	VSFT1֝cV�0M�� ��5�q� � ��EA_�  B8����E�� p�����ª�ÌB ��ME$�u4�����a{~&%��M���x[�p�30�$�xpTDINEND]H^8t�Or0U?��[J¨�S�ߏ���s5����Gy�	��,��������ߍ�REL�E �s/q�XOjFt�_ACTIV��~8��
 A �;}�<����RD�`��C!Y?BOX ����V�v��p2��>��190.0.���83����254�����`��� �q�r�obot�ę�   pHa�upc���u���p��r���ZA+BC�#�-,u�  �r�5X?Qc u�����/� 0//)/f/�Z;D�q���