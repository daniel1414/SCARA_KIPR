��   ?3�A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����MN_MCR_T�ABLE   �� $MACR�O_NAME %$PROG@�EPT_INDE�X  $OP�EN_IDaAS�SIGN_TYP�D  qk$M�ON_NO}PR?EV_SUBy a �$USER_WgORK���_L� �MS�DUMMY10   &�SOP_T � � $�EM�GO��RES;ET�MOT|�GHOLl��1�2�STAR PWDI8G9GAG�BGC�TPDSN�REL�&U�� �� �EST����SFSP�C���C�C&�NB��S)*$T8*$3%)4%)5%)�6%)7%)S�PN'STRz�"D�  ��$$CLr   �����!������ VIRTU�AL�/�!;LDU�IMT  �������$M�AXDRI� ���5�%.1 �%� � d%�Open ha�nd 1����%� a?�? �"  ��!�# �%CloseQ?d?�?�?�9}�7Relax�?��?)OOO�9�6L82 QO2O�OVO�3 �?�O�O
_�O�4O�O�Ol__�6�Fh_�_d_�_�[�3���_o�_ :o�_�_poomo�oUo go�o�o �o�o6H 3l-�Q�u ����2���h� ���;�M���ԏ���� ����.�ݏR�d��%� ��I���m������� *�ٟ�`����3�E� ��̯��𯟯��&�կ J����E���A���e� w�쿛�Ͽ�ѿ�X� �|�+�=ϲ�a����� �ϩ����B����x� '�u߮�]�o��ߓ�� ����>�P�;�t�#�5� ��Y���}������� :�����p����C�U� ������ ����6�� Zl-�Q�u ����2��h �;M���� ��./�R///M/ �/I/�/m//�/�/? �/�/?`??�?3?E? �?i?�?�?�?�?&O�? JO�?O�O/O}O�OeO wO�O�O_�O�OF_X_ C_|_+_=_�_a_�_�_ �_�_o�_Bo�_oxo 'o�oKo]o�o�o�o �o�o>�obt#5 �Y�}���� :���p����C�U� ʏ܏Ǐ �����6�� Z�	��U���Q�Ɵu� ������ �ϟ��h� ���;�M�¯q���� ����.�ݯR����� 7�����m������� ǿٿN�`�Kτ�3�E� ��i��ύϟ���&��� J���߀�/ߤ�S�e� ���ߛ�����F��� j�|�+�=��a���� �����	�B����x� '���K�]������� ����>��b#] �Y�}��( ��#p�CU �y� /��6/� Z/	//�/?/�/�/u/ �/�/�/ ?�/�/V?h? S?�?;?M?�?q?�?�? �?�?.O�?ROOO�O 7O�O[OmO�O�O�O_ �O�ON_�Or_�_3_E_ �_i_�_�_�_o�_o Jo�_o�o/o�oSoeo �o�o�o�o�oF�o j+e�a�� ���0���+�x� '���K�]�ҏ����� ��ɏ>��b��#��� G���Ο}������(� ן�^�p�[���C�U� ʯy�����6�� Z�	����?���c�u� ������ �Ͽ�V�� zό�;�M���q��ϕπ������R���
�Send Eve�ntU�5�SEN�DEVNT��3� �i��%	}�D�ata�ߘ�DATiA�߿���%}�?SysVar��OSYSVY��1�%Get��Z��GET����%�Request� Menu����R?EQMENU!�����?߀�;ߤ�_�� ����������F�� j+�O��� ��0��fx c�K]���� ��>/�b//#/�/ G/�/k/}/�/?�/(? �/�/^??�?�?C?U? �?y?�?�?�?$O�?!O ZO	OO�O?O�OcOuO �O�O�O _�O�OV__ z_)_;_u_�_q_�_�_ �_o�_@o�_o;o�o 7o�o[omo�o�o �o�oN�or!3� W������8� ��n���k���S�e� ڏ����������F��� j��+���O�ğs��� �����0�ߟ�f�� ����K�]�ү������ ��,�ۯ)�b��#��� G���k�}����(� ׿�^�ς�1�C�}� ��y��ϝϯ�$���H� ��	�Cߐ�?ߴ�c�u���$MACRO_�MAX:�������Ж��S�OPENBL �����՗��r�r�A���PDIgMSK�����Y�SUc�u�TPDSBEX  -�
q�U����n��� �