��   �A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����FSAC_LST�_T   8 �$CLNT_N�AME !$�IP_ADDRE�SSB $ACC�N _LVL  �$APPP  �  �$8 AO  ����z�����o VIRTU�ALw�'DEF�\ � � �����ENABLE� �����LIST 1 �~�  @!�$�����
[ .@�d���� �/�3//W/*/</ �/`/�/�/�/�/�/�/ �/??S?&?8?J?�? n?�?�?�?�?�?O�? �?OO"OsOFO�OjO|O �O�O�O�O_�O�O7_ _\_B_�_f_x_�_�_ �_�W