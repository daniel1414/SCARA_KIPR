��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
+GPCOUPLED1� $[PP_P�ROCES0 �� �1�!�U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $�,NO/PS_SPI_INDE���$DX�SCR�EEN_NAME� �SIG�Nj��&PK�_FI� 	$�THKY�PAN�E7  	$D�UMMY12� ��3�4�GRG�_STR1 � $TIT�$I��1&�$P�$�$5&6&U7&8&9'0'�'�%!'�%5'1�?'1I'1S'1]'2�h"GSBN_CF�G1  8 �$CNV_JNT�_* �DATA_�CMNT�!$F�LAGSL*CH�ECK��AT_�CELLSETU�P  P� H?OME_IO� �%:3MACRO�F2REPRO8�D�RUNCD�i2S�Mp5H UTOBA�CKU0 � }�	DEVIC#sTIh�$DFMD�ST�0B 3�$INTERVA�L�DISP_U�NIT��0_DO��6ERR�9FR_�Fa�INGRkES�!Y0Q_�3t4C_WA�4�12H�GW~0�$	Y $sDB� � COMq�W�MOJWH.�
 \�VE�1�$F �A�$O���D�B�CTMP1k_F�E2�G1_�3T�B�2GX_D�#� d $C�ARD_EXIS�T�$FSSB�_TYPitAHK�BD_S�B�1AG�N G� $SLOT_NUMZ�IQPREV��|G �1_EDIT1_ � h1G=�H0S?@f%$EyPY$OPc� �0LETE_�OKRUS�P_CRQ$�4�VA^Z0LACIwY1��R@Pk �1w@MENP$D�V�Q�P���A��nQL*OUyR ,lA�0V$1AB0~ OL]e=R"2CAM_;1� x�f$A�TTR�MP0AN�N�@�IMG_H�EIGHQ�cWI7DTH�VTC�U��0F_ASPE�CQ$M@EX�P;�@AX�f�C�FT X $�GR� � S!1�@B`NFLI�`t
�UIREs3�tGI�TCH~C�`N.0S&�d_L�`�C�"�`SEDkp;tL0J*DS�0>0�zra�!hp;�G0 � 
$WARNM'@f�p+P� �s�pNST� �CORN��1FL{TR�uTRAT@0�T�p  $ACC�1
� ����ORI	`!S<{RTfq0_S�B�qHG]I1 [ Tp4u3I8�TYVD+P*2 �`v@� 1,R*HD�cJ* ����2��3��4��5���6��7��8��9��qO�$ <�� #5x�s1v`O�_M�@�C t e0Ev�NG��ABA� �c��YQ������@����·�P�0����x�p�PyP�2� �����J�_R��BCb�J��2�JVP�CR��}@w��u�@nCP_}0OF� �2  @� RO_�����aIT8C��N'OM_�0�1åq38W ��T �#�d��@xP��J}EX��G�0� .��p�
�$TF`��C$MDM3��TO�3&@U=0^�� �H�2J�C1{�E͡� vE��uF�uF��0CPho@�a� 	P$@`�PU�3�f)�"��)�AX 1rDU�6�$AI�3BUFpV�o@�! |�plڶ�pPI��PZ�MY�Mf�̰i�}FZ�SIMQS� �/��A-�����kw' Tp{zM��P��B�FACTqbGPEW6��Ҡ��v���MCc� �$�}1JB�p;�}1DE�CGڙ�G�-�b�� ě0CHNS_wEMP��$GO����+P_��q3�p�@Pۤ��TC��{r��q0 �s��a�/�� �B���!�	���JR!0��SE�GFR��Iv �aR��TjpN%S+�PV!F�����ʹY��K��a1�)B���( 'j�Av�u�c t��aD�.0���*�LQ��D�SIZC������T��O�����aRSINF�����jq@��C��C����LW�8����x�CRCLuFCCCkpy�����N} ���bA�������d�*��DwIC��C���r���+ P��z�2EVT2�zFH_��Fp)Nt/�>�����H�1Q��!  ���Qx����U�kp��2 ��a��s�+����qRT!x @"�4�4u2��tAR��:�`CW�$LG�p���B�1�Pr�P�t�aA?@z�ϣ~0R�Ӳ�ME�`8�oC�RAs3�AZ����pb�OS�FC�b�`�`�FMp�� �0��ADIS+�aV%��b�z�@�pE$�pRp�cV�S�P���a+QMP5�`Y$8C��Me�pU��a�US" $=�TIT�1�S�SG1��#��8��DBPXWO�! T#��$SK���2o�DBTmTKRLS$l�Q0TQ���P`P�D�q�1LAY_CAL�1�R^0�o f7PL)A�Q�D�'a�73a�7���D�B!S%2?�PRj� 
*0���Sg& =�A$��S$ �*�L�9'�?H'�U�T(ODCS9)#ODENE��c*BO'Ӳ0RE�p�B+H �O�u�&$L�C'$@�3R��K2�LVO�s_D~!U�ROSbr�q�v�R����CRIG7GER�FPA�S��>6�ETURN�B�c�MR_}�TUbp\���@EWM$���cGN=`���BLA���TUܡ($P�')$P s�*hP3ab��C�TΣ@DO>����D�A���FGO_oAWAY�BMO"��a�!R�DCS�_P,<aIS t�� �� �s�S#�Q���Rw�cV��Q�w2�VW��'dNTV(��RV;����~��mgŃ��Jt��<@���SAFEڥ�f_S}V�bEXCLUT�:�� ONL���cqYfЀ�y�OTEu�HI_V} ��PP�LY_�q7�VRF�Y_b3� �Sj L�_G -h@0��_yО1� +�1�PSG�  .�rŐ1P NQ5�� _q���;P���Vby|rsvANNU�N<@�$�tIDX�UR�c[P� �y�qi X�z�v(2EF�PI<B/��$F�r�$А�OTQP�A $DUMMY��&����&���*0t�U0 7`  �HE�\����^r�cYRr SUFFI���Pa0�T�P)�5#�6#��1wMSW�U1 8���KEYI��4�TM`�A��ځ3QՆINݱ�v��1j P2 D���HOST�0! ��������������EM&����*0S�BL� UL��3 AZ�����)1T�@~S4 � $���USAMPa༥.������V I�@��$SUB����;@�c����3��SAV �����������`��vP$�@EC!	0YwN_B35 0��DI�t�PO\�M��#�$E�R_IB�� �ENC2_S��T6X��2������� �cG���0 S7�2��1��A����8  ��Ǜ��@�PK�Dk!uq��AV�ERҁ�����DSP�ܢPC?���2�6�\�����VALU��HE �M_�I�P(�ܣOPP� �5�TH��ͫ��SH` 4�.�FB�6d���~�� 5�SC?q����ET�9ȂF?ULL_DU���q�KP�ԝ�����OT��"T�PNOAUT5OS:�$YĪ�Z� ���X�C���h�CE26��V�L�� ;H *�h�L� �����$ P��wc�ě1�Ʃ1��@C��Ƨ��Ʋ���7�ɕ8��9��0����1���1��1	�1�1�#�10�1=�1J�2RX�2����2��2	�U2�2#�20�2=�U2J�3X�3��3�˪��3	�3�3#�3*0�3=�3J�4X�Jv�SE�2< <8�Z����I��e�$�}���FE5P?PT�= ,f��a? �P�?i��e�i�E�Pq�1azT>F�$TP$!?$VARI���n�UP21p? 7���TD��s��p��p��������BAC2@ T����$uP�*p��Þ0� IFIw� �0�P� � )PB"���0P�TAt ;`u�"�"pu STv t: �bt�@�l�6	sC2	>0���S����/bF��F?ORCEUPsr���FLUS�pHfN�n����bD_CM�PEv*IN_pt�e`�REM� F�a�a�0�TeʁKdN~�eEF1F�j�PINJa�wOVM�OVA��TROV��DT<	��DTMX,A ��P*��0M(xR#,�0�CL*_��u*ȫPr�{_XЉ_T��+X��PASaD% ��(װ�1`�&�_A@RQ�LIMGIT_�4�� M���CL�tˑRIV�W�*2EAR�I�OxPC�P���B��R�CMQP*�b =!GCLF�#�1�DY�8} �q�35T�%DG���0�5Iq�FSSt0��B PP��1�A��`_�1��8�11��E�C�13z K5 F�GRA��JgC��k�`W��ON��"EBUG�wctBx��C ��_E� D ���`��TERM�EyE�Eא�ORIS�@F�Eq��SM_��`���@G�EO��T�A�IH�Eb��UP>��I� -�Q���D|`�C|PE$S�EG#Z�0EL�eU�SE�PNFIz�LRT�kA,��DTF$sUF�`O�$\���a�P/���Wi@T���t �cNSTTP�AT��h��RPTH	JKa-�E
�65MR<p@&�WUw�&�Q�LQR<`<�Y�qSHFT��MQ|�Q�X_SHOR��*��F �@$�GM`H�u OVRq��q6`�I`4U� �aAGYLO���"J�Iu2�b��Q��oƸ�ERV ���a� 6j�WnP�R�~�E �e��E Rb1Pp�ASYM|�p�MQ#WJ`W�� E���Qy�b0�U7tnPI��Uw�/�ePo��`o�fgkORnPM�G@�SMTfJg�GR��aC�qPA|P��p|=��K � F�TOCFQ�P<9`N $OP@/�P�#��N �!O��ڐRE
�RdS�QOX����Re�R�U�N�%�a#e$PW�R0IM@��bR_p �L�=�mR LVB�H�_ADDR~$�H_LENG�RPǁ���T�R� SO�M H�S���~��������	�SEh!u���S:�MN�1N��p��F¹�OL��8�3�3�<=��ACROc�z �P$��[·a;�  ��OUP���r_�I���q�q1�ѭʓ�� ԙX!՘Y1՘t!՘	�0ԙлE"IO����DϗA�ߕ9�gO� $���p)_OFyFb�;�PRM_Ò}��HTTP_[��HjP (��OB�J�2��#$$�L�E�S���Q �s ���AB_�!�T���S�p;x L�V��KR32@�HIoTCOUBGE�LOہ磴!��@�0�"�G#�SS�ģHWD�SQjR��lpINCPU4BVISIO�����Ğ��
������	� �IWOLNS� 0�C$SL�r�@PUT_�$�@��PV0�ɱ)F�_AS�2T $AL  �� =a0U�@�9`dQٵ��䳊`H�Y#�]�6è��UO�3U `"�{�$�@5"M�5 Tƥ�R�P;@@��ǿ�T��µ�)��UJeV]���NE�fgJOG{W��DI�S��pK��� �3W� XХQVv��P;�C�TR�S:�FLAG�BB�LG�tX ��� ���aCLG_SIZ����d �����FD��I�اؓ� �׏ث@�֎����	� d 	��	��	�@	�% SCH_��R��ФaBg�Nє�Y���!E�2��p�J U�}�}��pL��|�DAU��EA�����t�▮�GH�r�p%�B�OOZh A<�f0IT2���@8�wREC�SCRB��=�D:�����MARG�<18��0��Ha�%�Sȣ$�W?��%���0�JGM��M�NCHz%�FNK�EY��K��PRGƾ�UF��g`��FW�D��HL	STP���V��mP������RES;	Hp��-�Cid@6r0�.0s��	U|����r�Xb��P�E���G��`PO�
.��M�FOCU�RwGEX,�TUI��	I��p�K|�V�� V����A`B���p��A`�Nu��SANAx%�FR��VAILy��CLP1uDCS_CHIyD�
��O�DX1�S� ��S�V�IGN��~�ӽ��\�T���_BWUFF�1[5�o`T�$��� ����RB�����A��\5��o`ܰ��c��pOS1�%2�%3�!t�|��0] � ܩ��qEU�����IDX�tP�bD�O� ��QV6ST|�R��YV�~@1 \$EO6CO;�{�^6q6���1^ L��K�[@`� 9`(��S���:������x��_ _ �o�p�Ð��� C�@C�p�` �� CLD�P|�uTRQLI���Ft
�4I"DFLG V�"@1VC�D)�VG�r�LDVE@DVEORG
�qiB_�g�H
�p�d�D�ta �M�P@Dr1DVES�pT4@�I��@TVRCLMC%T�O�O7Y���sMI��tb dy���!RQI�M�DS3TB�0 �VO�6�XAXr �X�\EXCES6��1vR)M_��qcg��RtPt�vR<��pd��V_A�Z��(k�_�X@K�te \����/�7$MBs�LI���c?REQUIR�b�x�l���hDEBU��*sQL�0M,�f�r=���`����%R�pMND���p�pgw�n�?�fsDC��IN�� ��p�,x' NV���K�sQ qPST�� h��LOCf�&RI���%EX�v�À�!�QsQODA�Q,�i X��ON���MF\����v9��2%��5�uk�0� ��FX�PIGG�� j �M��2!��h�3��4R �%?3�;�|�K�|�Z�G`E�D'ATA{'��E�U���b"���NZ"k t_ $MD��I��A)Ɔ ф��фH�p��`Ѕ�X�҃ANSAWe�ф�!'хD[��)�aO��P��l -�PCU��V�X@�uRR2��m D��a���Rd$CA�LI�P"�G�w�2N��RIN��z�<u�'NTEڰ�"nI����°r��ڰ_N��o@Õޒi�oT۔bp�7DIVmVDH�Pݐ:��q� $V��+sv1$��$Z�"���� �"f�_�e�r�H �$BEL�T>��1ACCEL�!������IRC���P��t�T31h��$PS�P'BL	` M�ʤ<C���������PATH������3ТZ��Q_�!U�2��8�R� C堌�_M=GP�$DDU���/�$FWh������q�����f�DE��P�PABNاROTSPEEH��!��4@�J��!��P��	`�$USE_���P���O�SY��g�Q �B�YNyPAO��OsFF��MOUR�3NG�O�OL�L�INC.��q��u��Rxn�PP�RENCS������Rȡ���TŠIN�'2IТ���`R�V�ES�{���23_UyPI���LOWL!A� �4@���D� @�R{`���0��5bCΐ���MOS4 LdMO����PWPERCH   �OV��b� �!m�@1�^T@1�s�� hP�`�� V5�'`ѡ��L���Ig�����UP�Ӛ���TR�Kv�#2AYLOA A��$a1�Т@�5�p40��RTI(a|�40MO����R$b�@N��T��w�L���"f��DUM2,�S_BCKLSH_CТ ��B�A�u�'�Y�������6�x���CLAL�z ���Ar�`�CH�K4@+5SH�RTY@S��}%�A��_:3N6�_UM(`n�C{��c�SCL��ʰLM?T_J1_LS��P������E�����p������SPC��0;���	��PCsѦ�!H�0�`Y�q�C3P�2sXTc�g�CN_��N��i��SH ���V	�*3�Ň�=Т�2AC� y�SH:3�� g��ƝA���s�4�ѡ���c�PAx�l�_	Pw�[�_5@��8�V�04AH�ZK�JGG"M���OG[��TORQU��ON.�Q靰`wbLҠᝰ�_W��1�_A��G��M��UI�I�IM�F�p��JPQ2(�A_�VC"��0�T,bS"1Y.�P8m/�R`%JRKY,�"��&PDBL_SMth�RM)p_DLG�RGRV��$G��$M��!H_ �#�:�COS;`�8LN � ;;\%B4G�=9M�=9 !y:g<-!�%Z60L�ƾ!MYD1�8$2TH|*=�9THET0�NK23M�BA�E0[CBFCBA�C�Q��R,B$:AG�:AFSqBG�XBEGTSaʱC��qW4&�Dxg3�Gv3$DUH� Ih�Aw�x�,b�F��,a9Q���v$NEd�AIF0Y�`R�E��$%��1A�5#U,W
581�LPH(eR��RS \%tSg5tSv5R�6�S(�Z�6%�VEXV:X7��]\VlZVy[V�[V��[V�[V�[V�YH�EX^Vdb\]�{hy[H��[H�[H�[H�[H*�YO6\OEXO�i[^UOlZOy[O�[O�[UO�[O�[O�6FR�'A�yg5�t8WSPBALANCE_�1��sLEo@H_�5S�P��X6�rg6�rv6PFULC�x��w��v5Ț1n}�UTOy_C�nT1T2G���2N*�z���g���@k���@ע����T���O����INSE9Gz�%�REV��%����DIF��1ol҇�1p�@OBȁ��#��MI��5��$?LCHWAR�����AB*y�$ME�CH0A�0>�D�Y�AX>�P��]�W(�<��q 
^������ROBV�CR�Ҡ�R='��MSK_�pj�_s P R�_��AR��H�Ҕ��1����ԲҐ����Ґ&�I�N���MTCO�M_CD n�t � P�ڀ��$N'ORE��9���(�ou 8�GR��I�SD�@ABJ�$XYZ_DA9Q<���DEBU��M���U�v �p$�C;OD�� ��o��J�j�$BUF�INDX԰MORœw $1�U��-��v�F���������Gܢx� � $SIMULX�����$����OBJE�p$�AD�JUSB�5�AY_	Io��Dc����G��_FIJ�=�T �������������Л�Հ�P��D�FRiI��׵T��RO���E��� ��OPWO� ɐy}0��SYSBU�PΠ$SOP���#��'�U&�ՀPRUN,�M�PA�DL�H�\!���_OU�!A����r�$��IMA�G��ϐ�@P��IM����IN� u£�?RGOVRḎ>�Ѐ�P����԰�@L�_:����m� RB�� �@M��E�DՠJ� ��NpMd.�������SL�p�ɐz x $OwVSL��SDI��DEXqk�i�=!{�$�Ѕ�V���N�Ѵ@{��Њӟךط�M�!=D�_SET�ɐ�{ @���g���R)I&���
��_4A���	���D�ׁ@��  �| HϑI�J�AT�US��$TRCp�@ǰˢD�BTMM�*7�Ij���4��#�\,�ɐ} DϐE~�k�A�`EۂBᏱ
��B�EXEH�Z�����{���~��АG�3UP���$����XNNm�=!p�L!p���PG&��!UB6�g��6�
�JMPWAI� PL��N�LO��j�F���#�$RCVFA�IL_C�j�Q�R ��Q�Z�M� 𣕠��޴0R_PL
�DB�TBm�j�BWD̓�A�UM���IGpe���m�� TNL� D����R���.�Ep��һ�!�DEFS}Py� � Lϐ�d�7 _: H�HUN!I��r�F ��R��^�V� _L��P@��	P�ȑ����F�����Ѐ��p��N�pKE)T�}�� P��ȑ�� hW�ARSI�ZE��l���S�@�OR
�FORM3AT3���COJ�����EMV�lUqX���D�PLI��~ȑ�  $#�P_SWI�-���AX����AL_ S��E A��B��,@C��Dj�$E6���uC_��	� � � ����qJ3�@����TWIA4�5�6��MOM������4�#�Be�AD�&��&�PU;@NR��J%�J%�DŔ�� A$PI�F �ޑ��$�%�#�%�# �%=D�&�+QD�DpсF����U���g�SPEED�`Gd*4f� 7167f���16g3�@8��O9��f�SAM��p맣417�3f�MOV���D�1ƀ�E�4�E$�17 1��42��� ����5n��Hm��3IN2Ln�39HUK0D�f�;J{HRD{K�KGA�MM�v�A�$G#ET��ȠL�D� �=
b�LIBR��]I��$HI��_��HP��bVE�XA^:P+VLW]XVO\:Y�|V+V�V����� �$PDCK��U�L�_�0�� � .B�m!E�W��T&��Yr �$I
�RS�D��&����(�LE�ޑ�Oh��)`��ѠH�ɐ��P��UR_SC�R��a^��S_SAVE_D�īe��NO�C����` �D��&�i��)�iap z{p���&Ex@� q��0�B���5G�2� +8!�;6��g8�w�ucs��1��DM{%� � ���!G����c�w���`ζ�qW�`��$��A0�N ��R�qM��&H�CLG�GM�aǒ�� � $PY�r�$Ww�+�NGt��w��u��u� �u��������@[�L�nX� O�mZp��GQ�Ŕ� pW�#�c�&�o�o#�5��_)�� | Wи�`������� �`�ޗɖ�EQ��E(g���b�/ ����P��PM��QU��0 � 8� Q�COUas�QTHHOL��QHY�SES�1[�UE�G��b� OM�  b�P4�U�UNI�.J� 2 O��)�� P�������a��ROG�j��2���O𤥥c�󠉠IwNFO(�� ��hث�
��1OI��� (`SLEQ�"6D�5D�ܦ����D$S𿠒��VPO�P�0j#3QEMPNU��Ύ�AUT�a��CO�PY�1�಼��`M"��N������CT��} �RGADJ(�e��X#�_$� ('��'�W%�P%�]`�'�:3�;�EX��Y%C��1@OՐ(�w� ��_NA�1!S���i����M?� � ��p��POR��Ì&��S�RV��)����DIT_p��� ��
�P�
�w�
�5�6�%7�8��1S�b��=���MC_Fe���pL�a�a�;�R q���/��җ#�0���k��� ,`FL�����`YN{���Mzp�C��PWR��������DELA4 �6Y�ADR��� �QSKIP{%�� �����OŀNeT�1�0*�P_�� ��I�`߂̐`��#`� 3`��n�kn�;�m�@H�m�U�m�b�m�98a��J2R.0��� m4� EX�@TQ� ���q����������jRDCx�� )���X��RF�E�@AY�_�X�DRGE7AR_�@IO�t=b�FLG���EP9C��UM_���?J2TH2N�# � 1� A�uG�@T�P �"����M��-�I���4�?�EF�11(�� yl!�ENAB� ��TPE2`{� 8 Wܠ�M�q�CL���R�w��2'��-?Qcu��3'������
�4'�'9K]\o� N5'��������6'�!/3/E/W/i/{/'7'��/�/�/��/�/�/�p8'��?-???Q?c?u?�SwMSK(�� /�t` E�aoMOTE���
���`/B`��q-CIOD�UQEI�0�p�qR� 9W\`��� /��� -�����ҿ���ՈB�$DSB_SIG!N'a�q����C��mE/S2323E���$��DEVICEUS�KC�r�rPARIT|!�AOPBIT�q���OWCONT�R���q�0�rCU�PM�sUXTAS�K�SNq��P�DTA�TU�p�RS�3`���u�e�_�pC���$FREEF�ROMS������GsETA`��UPD���AEb�CPTP����� !�8$US�A�����9h�{�ERcIO���`ՐRY�U�B_�`��P�QQf'WRK�?�<Dh�3f�h��6FRIEND<�qg�$UF�U��p`TOOLwfMY�d�$LENGT�H_VTߤFIR���cM�SE�@�iU�FINtrаAR�GIaF�AITI�i�gXF�i�fG2�WG1�� �Sr$wcPR��sau�O_�@�P��xQRE���SU�ءTC�N�=qyvG �G��]R���u��Q�A��hzhZUz��ZU�t���{P�T��X �P��L��TcH��hh�U�T�S%G��WX�)��r>�D���.��C�z�N��b��$�v 2!�!�-a' 3i1?h.`U21k2��31k3?j ���@i����6{��sL{��r$V��bV�e�V���vYr���O� [V{�@��hv3Ru�^p�ib��PS��E��$���c�5$A8й�PR)��u,��S���@��X�¯ 0p�v���P�N���A�!��P>p ��
�U�SzA� �\�RH��GA_�Š��Ny@SAXQ��Ag`L�a�g�p�THIC'ap��-����QTFE��|�m�IF_CH'c�p�I_����6D�G1@՘٤*��h��`��7_JF�PRW�I���RVATF��� �\�'�f`��)�D9O�e)�COUW�C��AXI�D�OFF{SEZ�TRIG�s z�,�)�#g���z��H����g�IGMAȞP�a\���ȸOR?G_UNEV#@Ͳ��SD���d� �$����GgROU[A�TOa��Q�DSP#�JO1GV�S8�_PV�3R�O���U�mpEVKE�P��IR?�_�=pML ���AP���E��8������SYSv��Bv��PG��BRKYr����b�\�������k�ADVQ�y�B�SOC�C@N�D?UMMY14��`�SV�DE_OP�1SSFSPD_O+VR���C~�N�&Q�OR\׶0N�P]ֱF��]�<�OV?�S!F��a����F���A�c�As�؁a�BLCH�DL�RECOV(M��P<�W�`M<��F?�RO1S�K�_a��_� @���`VE}Rt�$OFS�`3CV�@_bWDv� �`r���R��9�TR%Q�A�E_FDO>��MB_CM[A��B/�BLl�_¦�l��V�qDb�P����G���AM�Ú�yP��'��_M��>R��<HC4�8$CA2���|Ȱ��8$HBK�Q,��N�IO1e]�iAA�PPAQ�}�b����u��iB4�DVC_DB�c�񓡦B���D�A��1��'���3��^-�ATIO�@���FPM�UDc1�HFCABH�0bFs�p�p���Ea<�_BP��SUB'CPUk�I�S%��@ ����P�s�,���B~��$HW_C!���i��x�A'q\�l_$UNIT��l��AT}����I�CY{CL��NECA#���FLTR_2_�FIҤ�H)�FEaL�PU˲���_SCTosF_�F��
v��
FS�A���CH�AJa^���3R�RSD1�B ё�l�i@;_T��PRO ~�)PEM�0_���8�3� �<�*%�DI�P��RAIL�AC��rM��LOГc+�i���-���-'�PR��S{q�*��!C���@	&�F�UNC�³�RIN��pZ�+`? �$(QRA� mr 9��#��G���#WAR�:�BLuq�'4A;88�DA���!I835L�D�PA�A�q3h��!��q3TI���5�β��pRIA�Q�BAF� P�A���1��5��(T���EMJ�I1Q��DF_�`�ӨQ��L�Mt�FA�`HRDiYd�P�`RSoq�+`Q0EMULSE�`���E� �8��I���� p]a�$�Q$�Q ��,��� x���EGfP�AРAA1R�2)�09mb�E�50��AXE&�RO%B#�W�ac�_�M�CSY���Ae�VSW�WRذ�M12�� SCTR"Ņ�d�h�E�� 	CUq#��lqB�hP3�oV��)��OT��P� 	$�ARAYg��R_!�`	T��FI��j�$LI�NK�1w��Q�_�eS3�CU��RXYZQ��[��	co��Q)�R�X�PB!��"�Kd�
 � LcFI�eg3�D�9Ԫ$<�_�JN�"�e��SA�OP�_~T�[53�NqTBȜaNB�bC9��DU�Q�BV6r%TURN b���u�Q�!h�?�gFL)���B�@+pe�kZ73�I� 1�JnPKH�M��BV8r%p����c�ORQ& �!�#mX�C����������u��.�<��tOV	E�q��Mj�tC�zC��B�W�Fq� � ���� j�0���q w�P����	��q���0zC��5��!ERM��!�	v"E8P���#؄A ����id�%"�WP1MP1AX�bP1��&! �Q2�2!>�\A>���=� �`=�p=�ep=��p=� �@=�JQ=�@:�@J� @Z�@j�@z�@�� @��@��@��ב˙oDEBU�$�! �1(${�P��R�g� � CABP'N�[��sVְ� 
����Ϥ ��Ϥaڧ$aڧ�aڧ qڧeqڧ�qڧ�A�4p�`�2�RLcLABbb��u� ���1s �� �@ER�9P O� $8`� A�!��POB�FЉ�x�P����_MRA��_� d O0T<��\�ERR:���0T)Y�aIA�Vb`,�N��TOQ+�i�L�@H,�7R���� C�A_ � p�T�P��< _V1ْ.�V�2#c�2\�2k�ȱ���op�ˠȱu�$W���6�V�A���$�"�0,���6�Q��	�@HELL_C�FG�A� 5�e B_BAS��SqR��p�� �CQS��1�1��%�U22�32�42�52ڕ62�72�82��RaO �8��P,`NLzA��cAB��H �ACK��>�i���`�`G@ܩ��_PUr�CO,�@��OU��P0�`W!��3�7LTPX��_KAR���R�E��&@P W1�Q�UE� �p9CC�STOPI_AL �����Pq�Д���PGSEM���M�6��TY��SO��W�DI����}�L�1�_TM�MANR�Q��PEZV�$�KEYSWITCaHq8��CHE9OBEAT!�E�@�LE�$f�U4�F��5�K��O_HOuM�0O�#REF�p�PR�!)�AUP��Cr��Op�0ECOư|_1`_IOCM�d���5���g�@G� D�Q� U۲�{�Mw2Q��p�cFOsRC�3 �OM�@ � @����3�U[SP�@1(��$�@3�4�14¿NPX_AS�¼; 0�ADD' h��$SIZ�$�VAR2�D@TIPR���� Ah�а@J�� �� �BS���AC��%FRIF�a��Se�w	��N�F�@Џ@� x6�SI�TEFsj".esSGL}T�R7p�&A���#P~ST�MTJ�P�@;VByW�pSHOW��R��SV
@�D�w� �ԱA005p Ё "� '� '� 'T� '5)6)7)8)9)A)�@'@v 'V�	&r`'F( JP�()�P�(,)#`�(�F)p�(`)�p�(z)1��)1�)1�)1�)1��)1�)2)2)2�)2,)29)2F)2�S)2`)2m)2z)2��)2�)2�)2�)2��)2�)3)3)3�)3,)39)3F)3�S)3`)3m)3z)3��)3�)3�)3�)3��)3�)4uI4)4�)4,)49)4F)4�S)4`)4m)4z)4��)4�)4�)4�)4��)4�)5uI5)5�)5,)59)5F)5�S)5`)5m)5z)5��)5�)5�)5�)5��)5�)6uI6)6�)6,)69)6F)6�S)6`)6m)6z)6��)6�)6�)6�)6��)6�)7uI7)7�)7,)79)7F)7�S)7`)7m)7z)7��)7�)7�)7�)7j�)7�$�5�VPd��UPD��  ����)и�YSL}O��� � �`��Q��TA��8�����ALU���Ц�CUT��F��IgD_L��HI��IV$FILE_��?�+�$��S�A��� hҰk�E_BLCKh�x��>��D_CPU���  ��� �B�T���q�	��R �G�
PWll�� �LA1�S������RUN u������8�u�?����?�� �T?�A�CC��X ;-$f�LEN��s����f�����I�J�L�OW_AXIh�F)1f�,�2��M��	�G�_��I��Y�8�թGTORn�f��D��<ܣ\LACE��Y�pf�ٳY��_MA� p��3�	�3�TCV:�[�	�T�\�{�q�| ������	���J���ŉMĴ�J9�����	�r�2�Ц��������ΠJK�VKо�#���#�3�J0l8�'�JJ/�JJ7�AAL'�]�/�]�W�e4X�5��{�N1��P��M�I�ڤLӠ_��� b���� =`u�GROU�����Bd NFLIC���REQUIRE��EBU��b�Ŷ��2�c�	�a��� �� \A�PPR�C �ܠ
va�EN\�CLO��l�S_M`������y
a��� �P �MC6�{�����_M	GV��C�l��؎��5���BRK��NO�L�����R�_L!I�������J��P_��/��7��{È����6L�O�8���b�?��� ҍ�z��燡��PATH��������В���� $��ͰCN���CA �]���I�Ne�UC٠��%�C��UM.�Y��4��Ez�P���P�7��PAYLOA�J{2L��R_ANE���L����������R_F2LSHRC��LO��$���2�|��2�ACRL_� "� �����H�b��$H��CFLE�X_�`�Je�� :r���	�t������	�������F1 ���ïկ�����E'�9�K�]�o� ���������$��г �#(ؿ�����	TR'�X ˲�` H��%�&�8�J�\� `�i�W�{ńϖϨϺ����J��� � `������ʁ��ATl�ðELt �5j�J����JE��gCTR�TN"�F�6	�HAND_�VB�_����� $f F2�֋���SWy3`������ $$M���R �ӅH�ѕL��E:�F�A�������I��A(��݀��A��A	��@��۪���D��D	�P2��G	�qYST��yQ4��yQN�DY �Z� �ּD�E��)�����������H$� � �P T�]�f�o�x����}3>�� {@`���n�vf��o�ASYM$������Ͱ����_SH��#�=� '��dLHG�Y�k�}���J��G��gs]y��_VI/C�x�ӵpV_UNI���t�#��J��re�r���t ���t�ð	G�(H:j��#PX��2A�H��N��EB��3EN/@��DI	�W#�O���♀��� � �BI�aAK���� 吂��U��0`��n��� � ]AMEB\?0�g��aT��PTpi0��5�����AK�,p:�U�I�TKp��� $DUM�MY1�!$PS�_RF� i@$ڐ�͑LA��YP�V#��=�$GLB_T~@��ŕ5���`�8CAӁ� XI�	�֠�STȱ�SB}R��M21_Vɲ8$SV_ER��1O��#�CLߐ�EAuO炔��0O� � D Đ3OB���3LO�f��S�y�ÐS�p�1SYSS�ADR�1��5��TCH�@ � �,f L���W_NA�
����y5SR~>��l }J �J���F��B���G ���I���ID���D��� D���V�p�KYV���b u���ݻ������)�;Mt��XSCRE�i�W��E@�ST���F�}��a�Ǥ�w��0_�0AV�� TI�&����1�%������1���Z��O�PIS�1��~� �UEЄG� �񪠞�SG���1RSM_����U?NEXCEP�����S_ߑ��7��&�p9�T���COU\�ғ� 1֤�U�E��؂6�y�PR�OGM@FL�17$CU&�PO�>���UI_�H�� �� 8E��_H�E_������RY ?�0�����܇���OUS �� @��D�$B�UTT/�R����C�OLUM0��s�S�ERV�3��PAN�E�0V���TpG�EUA|�F��ʡ)�$HELP��bETER5�)��E��� Oq��30��;0��M`��0U`��]`��IN��-�ETpNp��0�131y� �i�;LN��� �0���9_����$H_�0TEX�3j�^�~$/RELV"D��~�Ԑ�b���Ms�?,@��p��4�򪑥#��USRVIEWV��� <���U"��]@NFI�0��FOsCUA���PRIx0�m��h� TRI}P��m�UN���Є� �`/��W�ARN����SRT+OL��&�Rs��O�cORNsRA�UW�vT�	���V�I�υ� =$��PATH����CACHV#LOG��LIM�r�Sx��BR'HOSTǢ�!���R|�OgBOTƣ#IM� ��Si@�0r��������VCPU_�AVAIL���EX�!�aN��} ~�`Ma�Ua�]a�����{0$BACKLAS� �!�$".W��  ��CT%s�@$TOOLǤ�$�_JMP�� ����$SS��v4ȁVSHIF`у�PB���Ǥ�Ї�Rk(�OSU�R�3W�RADI�$��_���%�м1��ぺ��$LU�q�$OUTPUT_3BM��IM���bp� }p���#TIL�''SCO�"�#C���$ N�&N�'N6N7N#8���u%=,B�2�P#�`Є�<���DJUrU��P�/WAIT���<���:%0NE~��Y�BOW� ��� $������SB�"ITPEo�NEC /,B@D(D�PJǐp�Rv hE(�#=@�0�	B�E/�M�KT���"`y�� An�!�OP�
wMAS��_DOآ�qT��D]����C���RDELAY��SJO�"X֡�c 'T�3��`� ��,l�y�Y_Ry�wR�#�ƢA�? �b`ZABC�� ���R��
 � �$$C�X����Q��Ȁ�P�PVIRT�_�PgABS�!��1 �U�� < �Q(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*��<�K�`�AXLM�TZK��c  ��]�INf�x�\�P#RE�Nk������LARMRECOV �Y�����@�F �U�P  dK��"� 4�F�T���w���������, 
#o�W��NGu k	 A   �,�`�PPLICu�?��U���H�andlingT�ool m� 
�V7.70P/3�6+��
��_S�Wr�F0����� 43�ˊ�yϋ��7DA7�철
�f��rm�NoKne����Oհ~�P�T����RAP_+�V��R�v�7�UTO�RX l����n�HGAPON��Pe� an�U' D ;1�� �и������T�n�� Q 1M�  ��������	7�H嵡]��R��R ��a�,�H��B�?HTTHKYV��R �+�=�O������3� ���!�?�E�W�i�{� ����������/�� ;ASew�� ���+�7 =Oas���� �'/�//3/9/K/ ]/o/�/�/�/�/�/#? �/�/?/?5?G?Y?k? }?�?�?�?�?O�?�? O+O1OCOUOgOyO�O �O�O�O_�O�O	_'_ -_?_Q_c_u_�_�_�_ �_o�_�_o#o)o;o Mo_oqo�o�o�o�o �o�o%7I[ m������`��!�[���TO��C�U�DO_CLE�AN��5Ի�NM  	�Կ��+��=�O���_DSPDgRYR��HIa��@����ϟ��� �)�;�M�_�q�������MAX@���[����׳�X�����҂�7�PLUGG�У��ӮS�PRCt�B�"�������O�}�^5�SEGF{�KY� k�v������Ͽ��8�=�p�LAP���� o�Y�k�}Ϗϡϳ��π��������1�v�T�OTALզ��v�U�SENU���� ����ߎ���RG_S�TRING 1~s�
�Ml��S3�
��_ITwEM1��  n3� �����"�4�F�X�j� |���������������0�B�I/�O SIGNAL���Tryou�t Mode���Inp��Simu�lated��O�ut��OVE�RR�� = 10�0��In cy�cl����Pro?g Abor�����~�Status���	Heartb�eat��MH �FaulAler%	U�CUgy������� ���۞����6H Zl~����� ��/ /2/D/V/h/z/�WORy��۲! &�/�/�/�/?"?4? F?X?j?|?�?�?�?�?��?�?�?OO0NPO��V@�+?OyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_8�_�_QBDEVYN�P mO�_!o3oEoWoio{o �o�o�o�o�o�o�o�/ASewPALT�q�/x� ���� �2�D�V� h�z�������ԏ�8��
��GRI���� B���j�|������� ğ֟�����0�B� T�f�x�������0�j�R�Z���� �2� D�V�h�z�������¿ Կ���
��.�@�R�ԯPREG�~���� dϲ����������� 0�B�T�f�xߊߜ߮����������X��$A�RG_� D ?	����9���  	]$X�	[M�]M���X�n�,�SBN_�CONFIG �9������C�II_SAVE � X����,�T�CELLSETU�P 9�%  ?OME_IOX�X�%MOV_H����REP�S�&�UTOBACK�����FRwA:\x� Z�,x���'`��xǣ��l�INI�px����l�MESSA�G������A���OD�E_D����#Ox�P2l�PAUSVA�!�9� ((O<������ ��(^L��p��ej@TSK  u����o��UPDT) ��d� ?WSM_CF���8���%�+!G�RP 2
5+ �L�B��A�#�XS�CRD/!15+ �������/�/ �/??(?�����/p? �?�?�?�?�?5?�?Y? O$O6OHOZOlO�?O|(�r�GROUN |S�CUP_NA��8�	r��F_E�D��15+
 ��%-BCKED�T-�O0�%_I_�� ����-r�_x��o�o�x���U2 r_/��_�_�R�o�iUp�_&o�_�_ED3o �_�o�_n_o�o9oKoED4�oro'�onpn�o�oED5^ �:n����ED6��o��npK���%�7�ED7�� ^����n�Z�ɏۏ�ED8J�*_��N_�m����m��ED9�[�ʟm7����#�CR_�����7�ٯD���ū�@�@N�O_DEL�O�BGE_UNUSE�O��DLAL_OUT� ��R�AWD_ABOR�𦾦A�ݰITR_RTNz����NONSi �����CAM_�PARAM 1�9�#
 8
S�ONY XC-5�6 234567w890H ��@���?��( АZ���y�u���\�HR5o�8������R57����Aff��\�L�^� Z��ߔ�o߸��ߥ���  ���$�6��Z�l�a��CE_RIA_I�(%;�F�!�{�x� ��_LaIS$�c%����@�<��F@�GP 1]Ż���O�K�]�o�.�C*  �����C1��9��@Ҧ�G���CP C]���d��l��s��R�������[��m��v��������� +C���& ��G���;�HEנONFI����@G_PRI 1Ż��T� ������ �CHKPAUS�w 1I� ,� BTfx���� ���//,/>/P/�b/t/�/O��x���8�!_MOR���� ��@B��%����% 	  �)?�/(??L?^;�"D����-=ֱ?99��3�@K�4��<�P������aÃ-8��?OO�J
 �?KO�'ưS����:Ov��i`��PDB� ��-+�)
mc:cpmidbg�O�d��C:�  .�P����Ep�O-_�C�  �  �KP�V�@�Oq_�<Z�  u�`��YU_�_=Y�,�/,�o�VXg�_o�]�,��S[f�_KoA�Mo�JDEF �ch�)�B:`buf.txtqo�Mro��0����'�	�A�ޙ1=L���jMC
�#�-,���>ss��$�-�r���Cz�  BHF3Cs7� C���C�M��F��iDP��E�~�WJI0D��tE�qaE�pIJ$�3H?HƷ��{�G�G��G�G���N[5�K~w)L��X�WI��O�fu7���4�),�,�.װ��,�,��@�u�K��x6�q�* RPd�D��n��pEWLI0E�X�EQ�E�JP F�E�F� G��}�F^F E�� �FB� H,- �Ge��H3Y���z�  >�33� ���|F  in6�|A@��5Y���<2��A�1WDq<#�
 �O+�)�Zj~�bRSMOFS����n6��iT1� D�E  �?DR 
��,�;�&�  x@�:��nTEST�b)o�8�R��!�/3��nvC+�A�WJq� �[��rq�C�pB�1 w�Cy�@T�6���T�FPROG� %ź��ů��I����𦶠喤KEY?_TBL  �6Q��!� �	
��� !"#$%�&'()*+,-�./01g�:;<=>?@ABC�`�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~��������������������������������������������������������������������������������������������������������������������������������������������L�CK�X	���ST�AT*��_AUT'O_D����G_��INDT_ENB�K��"R��i�[�T2<��\STOP���"�TRL��LETE�����_SCRE�EN "��kcsc��U��MMENU 1""�?  <���� |�WE[߅ߺ�V��߽� ������,���b�9� K�q��������� �����%�^�5�G��� k�}����������� ��H1~Ug� ������2	 AzQc��� ����.///d/ ;/M/�/q/�/�/�/�/ �/?�/?N?%?7?]? �?m??�?�?�?O�? �?OJO!O3O�OWi;�_MANUAL��ޞ�DBCO��RI�G�4�DBNUM��`�<q*�
�AP�XWORK 1#"�ޟ+_=_L�^_p_܂[�ATB_�� �$"��ipT�A_A�WAY�C
�GC�P *�=���V_A!L�@M��R�BY���4*��H_�` 1����_ , 
^7��6�Boo�f�PM��I�j��\@��cONT�IM��*���fi
�$cMOT�NEND�#dRECORD 1+"�qer9�Q�O�Oq =6��R{���Hx ��O�s(�:�L� ��������ʏ܏ � ���$���H���l� ~������Ɵ5��Y� � �2�D���h�ן�� ����¯ԯ�U�
�y� ���R�d�v������� ���?�����*ϙ� N�9�Gτϧ`�^�ϼ� ��=�������(ߗϩ� ^�p��ϔ�����9� K� ���!�H��l� ���ߢ��K�a���Y� �}��D�V�h���R�TOLERENC��TB�b�PL����@CS_CFG �,0k�gdM�C:\��L%04�d.CSVi��Pcl���cA CH z�Poo�n"W^m��c��RC_OUT -�[=`�o��?SGN .�Ur���#�05�-JUN-20 �13:34 �Q25-MAY��1:00 af P�X��n� �pa�m���PJP�{V�ERSION ��
V2.0�.11�kEFLO�GIC 1/�[ 	tH�P��P���PROG_E�NB�_r�ULS��g �V�_WRSTJN�`�Fr�T�EMO_OPT_�SL ?	�Uac
� 	R575��cO 74T)6U(7FU'50y(t"2U$�tH�/z2$TO  a>-�/{V_�`�EX�Gdu3P�ATH A�
A�\�/]?o?�kIC�T	aF�P00g|�Tdceg���1STBF_TTS�h�I�3U�Cda�6�@MAU ��b�MSW��10i�<(�l� ��2�Z!�mO |3bO�O�O�O�O�O�O�_tSBL_FA�UL� 3�_�cQG�PMSK��bTD�IA��4�=�d`���a1234?567890�Wc|6P�/�_�_�_�_o #o5oGoYoko}o�o�o@�o�o�o�o\SpPf_ *��OR*�?% �PBhz���� ���
��.�@�R�pd�v�H|��UMP4!fY )^��TRNB8KS��ĀPME�5Џ�Y_TEMP��Ç��3��D3����U�NI.��YN_B�RK 5����E�MGDI_STA�%�W�NC2_S_CR 6G��_ ����͟ߟ�f����`0�B���~�e�17�� ;������¯,R|�d�8G��a��� ����N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶�0 ������@$<��)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m���������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/��/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgO�/�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo�Oqo�o�o�o�o�o �o�o%7I[ m������ ��!�[oE�W�i�{� ������ÏՏ���� �/�A�S�e�w����������קETMODoE 197�v� '�� �W��RROR_PROoG %�%����X�'�TABLE  �A��������њRRSEV_N�UM ��  ����)�_A�UTO_ENB � #��j�_NON� :�
��_  *�F��F�%�F��F���+E�_�8q����HIS�h����_ALM 1];� ���F�F�+�� ��$�6��H�Zψ�_�%�  ��D����ېT�CP_VER �!�!F�j�$EX�TLOG_REQ栶����SIZ�����TOL  �h�Dz���A ��_BWD�5���a�	�_DIO� <7��	�h��k�STEPw߉�ې���OP_DO���4�(�FACTOR_Y_TUN��d���EATURE �=7�a���Handling�Tool 7� D�ER Eng�lish Dictionary=��7 (RAA� VisS� Ma�ster0�>�
�TEa�nalog� I/O7�>�p1�
a�uto S�oftware �Update�� �"`��matic Backup;�d
!��g�round Ed�its�  25L�Camer�a��F�� "Lo���ell��>�L,� P��ommj�syh�8�h600%�sco����uct%�ޡ�pane6� D�IFD�'�tyle select�;- `�Con��j�?onitor<�B��H��tr5�Rel�iab�� �(R-�Diagno�s���:�y�Dua�l Check �Safety U�IF��Enhan�ced Rob �Serv��q (�V�User� Fr���T_i�E�xt. DIO� ��fi�� Z�\�=end Errz��L��  pr�[r��C  P���E�NFCTN /Menu��v�����.fd� TP I�np�fac�  �
v�G��pl�k Exc	 g5t���High-Spe� Ski��  P�ar\�H��G mm�unic��onsn��\apur� �p���t\h8���conn��2�� !D�Incr�� strZ�i�<�M�-6< KAREL Cmd. L� �ua���8sRu�n-Ti4 EnvB=�(mqz m�+��]s��S/W=�"y��Licens�e��' a���o�gBook(Sy�o�m):��"MACROs,��/Offse��f����HG R��M1�?�MechSto?p Prot��do 5
$�Mie�Shif��9�B6SD�Mix ����7�y�Mode S�witch��MoT����.& �M�&���g' 65�ulti-T� �����Z�Pos��Regyio�  ! 7}Pr�t Funb�>�6iB/1��NCum ��dx�P`�|312  Adju�:�/2HSM7Z* yoY�i8tatu1�<�AD RDM�otN�scoveW� #��3��uest 86�7.�9oG � �SNPX b�����Z#LibrV�;�r't IE,� S$@��.�0�� �s in VCCM9��0�� ��!9��3��/I� 71�0< TMILIB��MJ0,@� �Acc�����C/2@�TP�TX"+QTeln� �Lq3�%|(PC�Unexce{pt motn��� �0�0,	7�\m72f�+4�f�K  h64aVS?P CSXC9�@�(P�U["3� RIN��We'50,�D��Rvr�	me�nS@� �QiP^ a�0��3fGrid��1play F �O`�fp@��vVM-��@A(B201 zf`2� ORD|��scii��loa-d3�41%�lJ�i�Guar�dP�mP���k7�b]aPa�t�& 0N"Cyc8��0ori���`{iC00Data�@qug�c�3[,`n�3FRLOAam�5�<�3HMI Der�2(�1oc644�0�PC�sePassCwo�aA)qp�1p����{-+PvenjCT����YELLOoW BO�I t�"wArcV0vis��x�%���Weld� �cial�$  k  �et�OpA �;�41\\�5a 2��a��po)@`@�a�T1���50.2H�T� @ xy�R:�82���`g�P��xp��� 12�AJPN� ARCPSU �PR\A�TEh0O�LwpSupg�fi�l5p�Q��^ l�c;ro�6 "T�`�3hELdx�!��SSwp�eetex^$ J�3�QSo�t� s7sag�% T�eB�P� ] !9M�Vir�t��39�V h	`s�tdpn6��roެ SHAD�pMO�VE TF MOS� O � Dg�et_var f�ails ��ߐ � � D��E��� �Hold Bus�tdCVIS UPDATE IR��CHMA 62�q��WELDT�@S� ) "���: oR741-�ou
��b��m BAC�KGROUND �EDIT Ò m�41�0REPTC�D CAN CR�ASH FRVR�TO�Cra.�s �2-D��r �0r�$FNO N�OT RE��RE{D � PCVl��JO�P QUIC�K�OP FLE_N .pc�c����TIMQV3 l�dm�PFPLN:9 燹 pl 2����FMD DEVI�CE ASSER�T WIT iC��sANġACC�ESS M �a:ŀo1Qui��<!:�C"�USBU@- �t & remo�v��<�2� SMB� NULApܡ��FsIXW��HIN͑�OL2�MO OP}Tt�PPOSTwp���D��- � �A�dd��ad. 	�i�o��$P:�Wu`.�$ѠO��IN��M���CP:fix �CPMO-046� issue�tJ�СO-|�2�130����SET VARIABLESΐ��$O�3D m�"view da`PW�ea�80b. of/ FD ��u)��?x OS-1�p� �h s v�D�5tv��s ��lo ��(� WAx��"3 ?CNT0 T�S$3Im�Z#ca��PSPOT:Wh�p܎�s�STY܄At��pt�do G�ET_l���VMG�R LO�0REA�pC��M`P�@ �Y��0�ELECT���L��ING IOMPR N���Rɰ�̐sPROGRA�M�RIPE:S�TARTU�@AI�N-��D��QASC�II�d�OF L����!`PPTTB:� N��MLKdme��4��:�moW�a3ll��R� Nu�Qr� Ang���`Yd��tho�n[� ch >`ܐ�r �R2toun�H85>@�iRCalA�"OSign�0�pI,A��Thresh1[23�#.c�Hڰ� : MSG_P�єper �ࠡ��=A�zero5P� �A�  J�!O�Im�r � 2D�0rc �imm�`SOME�s�ON������0SREG:�^5�� LB A9�KA7NJIH�no��`9c	��n dq��� -1o��INI�SITALIZAcTI��we�,�0= dr\  f��a|P���minim90rec 1lc0��:?!blem��r�o��L�<3a i� Q09 ��b�d�w-�q ݡ�0�w uHQ�m@se�4SY�M`��s���QЧ 090��Wlu� E;BRe���jձ4�1���m ���Par�r@ G��Box fo T�ME�ːRWRId<���SY��\k���F/�up��de-/rela2Qd��#�5�betwe�pI�ND��GigE osnap�us5��spo V�TP�D��DOs�ġHANDL �`�Q�i��D��n�0 f.v����Boperawbil�` tmCQN��: H5@�`l��L�
! ��m@}ph�s UIFL�PO>�FA����ΑwV7.��CGT��pi�AsM�5pj�)@�U��ine-Re�markO@0 R�M-�$ÔPATH� SA̐LOOS����v�`fig�G�LA  �0%���p̗�J� ki q�thser�A� Tr�`�in�DW����2�7�� X�е���8`Mn;� C� ��:  �6�d� y* it �35\k�Pay΃a[2]_�D1:� g�s> dow�D2	SDISp�1�E�MCHK EXC�E ֠�$MF +$  ��h�"�P�����B0 ce1ȢF��me�� �c� �!?��bP�� BUYG��yB
�@DŠ�PET��V0�0�T9�3X�XPANSI�)�DIG��O � H5�P�CCR�G ENCCEM�ENT`�Mm�K �1A�H GUNC'HG OA�1Tڐ����Sg\d���1�0ORYLEAK𯱄���LC W_RDN R��O�`sj5`PO�SPEް�CG�V ont��VM����W��@`GRI,@A�7��� ��PMC ETH̿0i�SUذ>� H�57�P0PENS�!�N���ː RE; (i�ROW<�³�RMV ADD c II�=p��DC^ ~q�T3 ALAӀ� ��m��VGN EARLY>���f �n� ��衸E�ALA�Y7u�СPDg�ˀHz1SS8�OUCH��D��Fh�����PCD�ERROR*PDE���� WRO��CU�RS�PٰIp@N �gҰ�?Q-158rKwa���SR �rġU3��\aptp��@T�RF@�R�\`�UB�U �`��#R�B�0SY RUN�N���`10�ఱBoRKCT@qROq�0Ԁ���CDAX��D<jj�EISSUcހ�\��D��TSI�aK��tXM�IPSAF�ETY CDECK "M6���d� ��[`S U�)��4}P@Q�TWD��E�'QIN=V��D ZO�����a�sb_aBDUALP@|�'QòF��E�4�l�6��P`NDE�X F�P�U���SU�F�rPk�Lbѳ�RRVO117 Ay��T��챤 ��FAL>�BTP247����P?q�EHIG�PC�C n��0�ESNP�X*PMM�Q ��)!SQ�"V��8T�bDC��BDETEC��d1s!Sˀ�BRU/b6x3���s� 02"�tH�s�'�!h� Z�T�7�pS��"e���߆���,����߉ـ�0�
�ա��ق�cscr��ـ �dctrl�d.؁���f$ّ��!���fـ*���878��-�% ^��� rm��
�Q��R��78�RI0ـA�̑ (��~�@�Q.����ao�ـ\���a:P���a��I��t�a 3 "K:�����<�#�o��tp؁ ?"PLCF"E!�<ـ�plcf���8ـ-���mai�ـ�N���ovc���ـt �/�ـ������􁢐�r674��Sha?pe Genwـ�I��R,���ـT�іV� (5�ـ��II���� �+��ـ�l���sga 4P�3 4j�I�r6ـŲ�5=�5ѺI���et-s6� " PC���{nga�GCREѿp|�5��@�DATj���5ŝ�t.!��5��a񯜳A�gtpa�db���Y�tput�������ñ��2�ـ��5Ĺ�����sl��q� 7�hex�y��4�����2�ke1yy�ـ"�pm����f��us9ߜ�gcـ ����+�H�a��j921��pl.Colly󔱾�r�bВN��ڕr� ({�ـip���r��'����8�7=�7���t�p�� "TCLSxj�|���clsk��tD���s�kck�� �)�U������r�H����71a�- KA�REL Use {Sp�PFCTNj��7��a�a��� ( ��ѡ�� �ـ��ٹ��6�8=�8"   ��ـ 0S��(V�   3lm� 6�99�~ �F�)vmcclmf�CLMl��`��60fvet���LM:�̙��sp]��mc_mot���ـ0y���suX���60���joi�T�J��_log8H��trc��ve%�� ������g�finder���Center qFb!��M�520��ؙ�g��  (m)r,���fi��1�� a#z�� �ـJ��$�tq� "FND�R����$etgu;id@�UID�ـ�
?1��E7�q1nufl�6 �ـ>_z#ѯ7A�x���(�2#���$fnd�r����c$��tcp<S$]�CP M� H��3ـ517��g�38�vC�gD�*Y= �F| Ց� ^ ���CtmgA4�P��O�C G1ՑO7�Y��8�ECtm �?�Wـe�?�C�Rex�ے��p�Z��ڔXprm؁��_�D�_vars �_Z$M���Vh@����`�gG��ma�w�G�roup�@sk Exchang{@�ـÖMASK H�5�H593 H�a�H5���`6�`5�8�a9�a8�B�a4q2���b(�o#
Ak�/�غ`hp8�0Y�0/_цt�qTASK Y_�r��pz�h�Z��m@��������SDisplayIm��Qv{Gـʑ8�OJq(P%���@a���aϘ� ـlqvl "DQVL�t���q�����Ϧ�y������1avrdq8֏4ᩅsim���0F��st��o��d���������v�0Z樁����"v�Easy �Normal U?til(in4�|+11 J553��a�c���(���0��)�M�<�O�<� k98�6TA8��#�4�� "NOR�
��1�_���|�su��.�������7���a!g�y! mOenuu��g#M������R577� 9{0 ̒J989��49�L�A0�(�ity�E�A�,�P�mL&��mh8��"8 2 ��܄����C8_S�շ�n "MHMN�r%.Ը%���ͯ�s@����i�Ը-at�Ѐ�_�������ֶ��tm�?мz�1����Qđ2�Ͽ�z�3zos�ogdst��
�mn�O��ensu�Lm���hRaL�߃��?huserp�a����c~���Ը5�ɯx�����oper��|�XԸdetbo`� �~ ��LUA���������dspweAb���+�X���u<1��101W�הּ�12N�A�e�30A#0�D���4N�;2e�5���|����"��Cal xN�0�O��Z��0�O�$��S%j{�u���� 0S�}���u�mp��\bbk9�68�!68�!��b\�eq969�9��%��F0b�� "B�BOX�ۍ�sc�hed����se�tu~Xk��� ff H)�0�eq)��0�col(�1bcxc��8�li�� ��aI���W!i�e@�m�rof$TP E�B!TA&@ry|M42�7�*l!(T\�Q!RecX"H
�qz�?$it�%�?#сk971��!71�{�F�$parecjo��A���?'����Xrai=l�@nage��~@�]��D2E� [0 (?:H͒V|x@1ipMa����3�p�!4�"4��u��3paxrm?r "XRM$��3�rf�Ͼß1�1�ꫝ0�yturbs�p'G#��^@ �0195: ��625t/~A ��\BH�'ZDiy!:k�E�6�"A���H� ��7��P�.�E!pd "TSPD�}<�T�GtsglD���kY��O�CiCsRct%���HvrvQ����K�P,��A  cq#-a21��Y@AAVM l�r-b0 �fdE`�TUP him �(J545 �l) �i`616 �V2VCAM �.CLIO �Y10k 5W` {(F�`MSC ����bPs�STY9L�Sua28 kr�`�NRE I��`SC�HgRpDCS�U tpsh ?ORSR �ua�04�EIO�CW`\fx�`54�2 LEX"�`E�SET��iay`0s�hi`7y`"RM'ASK�b7o�-`�OCO[�x�a7p3PSv q`t7p0kv6U`�xv39_v�xLCH�RvOPLG�w03�;uMHCR3MpCе`YaP`�p6�.f�ia54; #�MpDSW�`588�ip1��a37 88 (%Dr0c�5r4���r'7 qj5r5�5r�^v�p5�"9P�RST VRFRDMC�S�a��-`�930 ��`NB�A  g1�`HLBo 3 (�aSM��� Con�`SPV3C Lia20�#-`�TCP aram�\TMIL �r�PACC�TP�TX �p�`TE�LN 96�0�r9^/uUECK�1r�`UFRM etL΁aOR ���`IP�LKeCSXC�pj��qCVVF l �F7�HTTP satrbZ0zcpCGy��8�AIGUI��p7 ��PGS T�ool�`H863 dj��qM�Oq�3
vJ684c�\�$���sق�s'�1�ےs�a96 TF;ADȑ651�Cq�53 � oo�b1B�44r-�k�r9��VAT��J775� �R�6uAWS�Mے�`CTOP ��q�`old��a8m0;!diy�XY�Y�0 e��i`885 '��`L�`u"�`�� 7H�`LCMxKP��pTSS J�%�
�W�CPE �\dis�`FVR�C m��NL�Uo002 
�en%�O6 65Jr'�7[�U0�po�ࠠK����t� I�4 URI�5��&�U022 n�se�{�3 APSFI�`{�4�2�`L-���alOP��1C��33O�͐tpts�D`U040g�43��ٲ4�۰j� "Csw%�1`b	�4�C�	�5 ��wx�57��eU061��S�6.ұrob9�5g�i���68����!!��7��w�7�Ё�%���"/rkey��3w��A4?ǽ���T���8'�w089�U09��d�P��9:���2 &�Ul �9&�l��9B��VrU15�P�M� s	lA �3#�}��ũ1q�0v4�7��1�08 	�eэphHc ��s�1�q�4+�Q1����A�5/�tx�)1����1]pu�Qф��t�1�����`��3����6��1!p �`��о�- W8�147 ase C�xU`sB�1 82���1�4�8 (W;ai��59 ��a'U166�W�1�W��4� j U�6�#U�7�3U�8�3ѱ��B��y1{��2 act�~��6 "MCR@ِ҄4�1������9{67ǑU193�3���6��2Y�sP��2A��21��as�F���<�2-���E�'2 wF���55�(���� ��cر5)�w@���q��p����qf�� L��$������q4d��!2g�8q��8�51�""@]�}�q��< b������B]�� f��; `�̑ � 8 16 (ݰ�BA� �AAҰ�]���g �:�!��`8 bb�fo=� t� j�� 7? \� ]��� �2 k_kv��74 &!����fW0H5��57&��579 h� L8�2 %"��4K 3��5����5��x1��594 U2N19 7,-�6�pz��6i�\tchH�6ur% �4S3� 90� h�&��\j670��q ���r!tD�4���&�t�sg�lIc�S�FrE�H���#F�����hk $�� sC�� ���"F�L��dflar��� �� �@��fu!l%�gvPva����sA�����"D��3��!creex���!�%�!`�%�,���6j6�=s�!prs.�!�% �!5�hA�P 5�fsgn��/�/�,at<D�AD���q|s`R svsch`@�Q!Servo Sμ!uleoCA5SVS�!44���F���1 (�0Ached�0,1�EA၍�� �2Q��0��^�r0h�U)1BBc��� %P5)Q1�V-#�3�1�css "ACS �WVY88"gA�`8!�/�0��@e�Ҿ#M��C��3�torchmܤ0�- TQMa��1�1M%'�9 J5^lA598 א1�!7)P8<P(1̢A�pء%R1Qte,�!�)E A5E`ASv�� �mLC6ARC_�k 1�4q� �V,�Ht!tc�A耥Q8�4��R F1 57T!2�SEPBPQ8f-!�RtmkQ!p@c60X��/�PRC8S��Q#�S�) P�2a9�6xAn`X�D.<bH5��1�U�}E� T�Qf #` aQ!<���F!�T!!a4�3FcRO�Ttm �R!av`58�_�WP��MA$q�E8��>rp�in_���o�@e`AcB�rr�)u�!�U�etd�ѧ�U>�Qoveto�#$,��S�mmonit�r42�=�Q�c�st,"M_va�P47M��V�0�! 5�q����ameQ!Ɂrol��A��43$Q0 � Sp��1�01$P2y5�AKR  ��� 0S�(V��Ɂ)xj818\nl`mD��zN��r�MPTP"�O��qmocol�]/
� Y1�4Xa�@��2�0i��53(1��Touc�h�!sؠ�2%qD2J5 !IU�٠��= b�0n��A��]�vP��`�z�EOWJ�th�Kwc���{�et{th8!THSRX���m�t�o "P�GIOsRd�'z�wk� "WK1�aL&�MH�PH54�5�Q5�o��m`A��q@!7z@6���18�a�P�Mor��tsn�@T �A�o�c���"���
��m�uA��T��p���T?�|�m4�TM�!2�54�>��� �m9�w�f��S�3�G�qor�3���"641���8ⱐQ!A�,HE!pRU <��m�Re�h-g "S�VGN_��(copy "COTA��U(���r#j0 "FSG@��_�eh��f�@�wA�SWwjRbY=sgatu���!�;Bv�tp�ATPD7��9 a79s����sg8!��GAT�&o<Rc9  �Ħ�1�t2`%1��&��1�bpv�1��& �1��B �1� 6�1�chr��1�|v�1��sm��1�v���gtdmenps1�(v�0!1��mkpdt��r1��]A1��pd���1�$&�1��m?vbkup.1��6x�A��mkun���G�pr���mklh1�e�P�s1�ni��<0&1�ldvr���glg�t�1��&����#�auth�.p �&��1�����) sud�1�7� 1�G��1��\1�g b2 �p�w 1�6O�Ł�4� 1�Ђ ?  946"1�����1�t\paic\p4k9471��wc��1�ict3as-�Mpa�cck0m	�	'gen!1� w�l��Q� st1fq��q�wb����������vri /�4�^��B1�D<��Pflow�@���Ac0ow�3<R�50?���Q�TR�  (A0e T�)B�Ԗ�cud!�w�1��fz�ac�$046 a0� =�f�+paRa0���!1�355Ţ1���F�ѡ�)a%��;:aOfcald� �&��0����%�f�m�:�"�#�4�`��'a�`"�3U���$�B1�!? track���@�aine/Rai�l TrP��{(699�/�@ (L !iE YB�ʔ_VB!BuŤ�a YB38P�4A8'7�	�F2��4�P�/�C�B1�3Ţ3�/��IUal��1�NT`����VA��zQin�p8�?0HVaen0�? DXWApuA�YqBzQtstd�0U�@1GW  ��]�j�VD���E&���VH@���open�ers^CO�`�AD#ev/w'~6�F8���񭁶��bA�aes �#1�]�ג�d���0�m�d1�k9�@7��6��#1��/b�epwaop`aOPN�Wpj�`��Krcel}?�Exg���Y`5Dv��tscx?t��a�sz Fuvrop /�Dw�nDh��bAr 5��QB�g�dk�j!�� Pumpv$Aᛑ��/�1�a;��M ��T�q�i���tx4U�1� 0S���O \mhplu�g�gr7Gh���uX|bZ#��ioh#C{p���v(�ALIO1�1��@7��93�Q5�1�91�����4�� �ST�
R�t�J9s89��/RLSE�g�1�@Cd�(M�1�/O�'�Q�)�D��G1a zq�H155'?���zq�tcmio���MIO�$�t}c�q"CL01�U�QcP�|�io��u~0%�l9�zp��Dv�1o���Q�tzt����dtz5I$��xV%�rh#Inte�Q.�� Co~Po�qv�RP1�hd�B554# (l�oBv�,�Q�H��Tcipc�oo�ڱp5�A�(
���������"7`���aڰd�QCD�W�	�����8��ڱ�rcnd(�_׳1p�a�ײ@������S��a���O�2kz�rp�crt�ᱯ�pٱd Ec��S d�\���u�xE!߳vr2k�p�E A�-�x�_B\"� c3hoO�l"uC��Y 1খ630@ᗷ�@ �� �ӿ�q��ԑ�G�TX�? �Е1ch�p "��XOh:�3��&�"5x!E��\p3 ���P��j�d �11�$h��Plo0���ұ�ch��3��s1��a�01���#Ar��0� !oCB��spq[Jm:�k�7�)�vr�Ҿ���a!�X%-J�FRAJ�W;atpqrnev'�����fQ��D5�`��KrboT ,�$��@PG�[!�sm�ICSP\QQP5y�x�!QP����j�H51z�93QP7y�6������2��5��R6QP����NPR�`(P@aam S`u�b��ĉ>a4tpprg�p�B�	�Z�qratk9�32(q v��sc "iC��~�atpr�_�qqz��;F�LGdsblf�lt{�ёsabl�e Fau`��C�Pav�aQ��`aDSOB (Dt$�t�d �A����QPh"�E1��`f$*��3[S� A�"tdj  "PaV�Ohf$�1sbj!��1�"\:1gc��.�f%�du��550^CAdju�st Point�b��J/��-�0�4��a昐A��j�O�N0\sg�4��w�1�\ada��"AD�J�M�j0�ets{ham�SHAP0���XDjpo �e��G �a��UGQPG'.��1:��k@ab5�J�KAR�`�iagnost�i��!�a��66 �J�C��a=P(QL��Q&T�o�fkrldeP@���	 ��SQ�$�)�3/ρ[pp��ODBG2t�!O �U@�Rѯ#��V��F( �Ѱ�S7��Q�ip{�M��ipper O�p��Pq����78 (MH Gw�1Rlb k_�fTcBQ��0&�d038<B8t��E��c�9_9t��Tc��k����8$q�Sd rnpVǁ��Qd����6Tea�=���r M�at.Handl�v �an`W�� MPCLGv�A_�p�q(�s є�f����g��b� �a���f������ >@$w����Dw��EI  d���uu�m���fhnd "F��?  ������#� ��p��>��(Pa�0To@�$V�!!�3#p��a>��{�^Q�k925��26�Hq�3�{�p����2	Ÿ��y���gse>0GAS�qďėPR��T��0��a���tp����{�dmon_�q�Ŗf�ans���vr�� {�=�����ͪ�<y��w�sl� � pen���D��Y�WA��823X�Q
�G�0!'� &P��8QqIQ�GQ �\sl��!q�� v���������֐�_��`����"SEDGpiOٳaQ�tdg�@T�AF8�F���BN��� ÑQm�7���ڱA��g;Ж�Q�����q�S�'ileg�y�e���π��9�F'QQ�LaQQj�517So�3-[J@V�?�'�#4A�49GA�WL�aw {�nao�Qfԫo�H17D��#a�����0t��  >��LANG j��A5��5�5� g�ad5��C5�TC5�jp .5�ce���5�ib=�5��#5���p�a5��C5�WҸ�j5�39.f5�]QRu~5� Env
5�5S��K�3y ��J9$5�.� �;��G5�2D25�JS���p(K}�n-TiAm��"���"��3H��������\kl5�U�TIL"�����r "QMG��,q5�8C5��1 "5�ړ�5�s5�\kcmn���+��r5���ut|M�_�lread��ex����"��\"��l$"��135�rt[! -5�tuva���`_��5� �`C1V����\p ����Bp9tboxx��_qcycs}�kRBTvveriOPTNv��l��e��K����hg/�ag�p.v1$�"1$pt�litDPN�D�BPm$dn#te\cym$8$o"��#mnu3�/�/�/�.�5�/�/m$��UP?DT ite��.3 swto95]�-4oolBD5wb95���-4FR-4Y�� /2gr�d�-4��-4�b-4��w -4B-4.3��-4�@-4'�-4�.3B0l� /2bx "�5�Q5I.3tl�7��AE�#/2r l\�6�@O��-4 :4ColD5eMa-4+�C�5K�-4W��Q5ml�-4Chan�g95}�95�qQ5rcAmdE�b�OZ�`6�5,r�7�6��7�5&r_&+]22=_O]2� c_du_3U4<_N^57�_<�_1UCCFM�Ey�>�_accdau59#�6cAEX`�/2|�D a��4|aO/Jm�a�5 �-4@�4�aAOSJ	Q �e�o�oY��-40��ZDQ-4sk��?
�@rtet�q-4\$�3<�q�eunc.-4�8�4�q�5sub�5��85E�q�5cce�@o�Rf^opm4E�o�fv �7�o�eT �c�o�nt$ 
Pte;�q �@�f�\��k��6;�-4�� -4K�D��z<h!-4xmov�b��q�et���f�"�tgeobdt.���ƥ�etu� ɐ��$ɐ��tɐٓxߟ�9z��var'��sxy&��pclJ��cɐ��ɐ�eɐg�ripsu����u�ti�����infCpo��ܯ�ɐ������\����ɐ����8�p��n��ɐ%�ɐZ�mT���ɐԶ��\�ogġ�Ʊ�%�p��\�palp�����s ����ɐݵ��Ŵ�����p�p����pkag�d�%�7�lclay Y�k�A�ɐ��dɐ5�p�������B��|��|�������q����rsdmͿ��rinT�-�?�sO�Q�c�̿޼1s���ߧ�tv�ߧ�qh���stn[`���tX01ɐ)�D0ɐ� �Tul4�q���g�26Ϥ�upd����vr����נ�1}�3�נ��ϵ�i3l3C�U�l4����T�5e�w�s ߘ�֠�߻�wcm�(���xferϪ�tl�k2pp��cosnv�朗cnvݑ���5�ag, y�l#ct���n�p��nit0���d��Ǽ(��  �ɐ �0S�(V�lU9al �pm�Wse��2���� V�C��(�z���A�0�|�m����&$��޷'#ro��T/f(&���p1�mI��,�� $�+���/�)G�?@�+�� �L�ɰm � ��P?b6D�4rg� ����������?�9 �� O�7����� �>�/�T�a�8/�C �����E��b,֡)?�*��nq?_9l�-!H��  �HA� |�p�QU1 p! O���P; ��S 	�Q�R�@t�`  �?��ɐ8?� �M�.Oreg.ԃnO��o99 �� ����$FEA�T_INDEX � �S ����P�5`ILE�COMP >����ba�Pa�RUcSETUPo2 ?belb?�  N �aUc�_AP2BCK �1@bi  �q)�R�o�o  %�o�o�Pe`�o)oe�o U�oy��>� b�	��-��Q�c� ��������L��p� ����;�ʏ_�� ��$���H�ݟ�~�� ��7�I�؟m����� � ��ǯV��z��!��� E�ԯi�{�
���.�ÿ տd�����Ϭ�*�S� �w�ϛϭ�<���`� ��ߖ�+ߺ�O�a��� ��ߩ�8߶���n�� ��'�9���]��߁�� "��F�����|���� 5���B�k������� ��T���x���C ��gy�,�P���qi�`P�o }2�`*.VR�H� *Kq�w��2PC��� �FR6:���/�T@`@/R/��=/|,C`/�/�*#.F5�/�	��/� <�/$?�+STM� D2M?X.�E?�=�� iPenda�nt Panel�?�+Hz?�?j7�?�?8?-O�*GIF7OaO�l5MO
OO�O�*JPG�O�Ol5�O�O�O5_��
ARGNAMOE.DT?_�o0\S__� �T�_@_	PANEL1�_�_%o0�_o�?�?�_2orog`oo/o�o�Z3�o�og�o�o�oH�Z4zgh�%7�KUTPEI?NS.XML�o_�:\���qCus�tom Tool�bar(��PA?SSWORD��?FRS:\k�*�� %Passw�ord Config��������+� �O�ޏs������8� ͟ߟn����'���ȟ ]�쟁��z���F�ۯ j������5�įY�k� �������B�T��x� Ϝ��C�ҿg����� ��,���P����φ�� ��?�����u�ߙ�(� ����^��߂��)�� M���q����6��� Z�l����%����[� ��������D���h� ����3��W���� ��@��v �/A�e��� *�N�r�/� =/�6/s//�/&/�/ �/\/�/�/?'?�/K? �/o?�/?�?4?�?X? �?�?�?#O�?GOYO�? }OO�O�OBO�OfO�O �O�O1_�OU_�ON_�_ _�_>_�_�_t_	o�_ -o?o�_co�_�oo(o �oLo�opo�o�o; �o_q �$�� Z�~���I�� m��f���2�ǏV�� ����!���E�W��{� 
���.�@�՟d����� �/���S��w����୯<�ѯ�Ơ�$F�ILE_DGBCK 1@��ʠ��� �( �)
SUMMARY.DG篞��MD:�[����Diag S?ummary\�i��
CONSLOG�Q�4�F���߿n�C�onsole l�og�h�G�ME?MCHECKտ���J�c��Memory DatadϾl�� {)O�HADOWY�>�P����t�Shadow� Changes���£-��)	FTPҿ?���C�n����mment �TBDl�l�0<��)ETHERNETaߑ�"�����n��Etherne�t ��figuration��s�V�?DCSVRF`�F߸X�q�t�%6� �verify a�llt�£1p�1�DIFFi�O�a����u�%��diCff���"�6�1��8����{� ������	9�CHGD E�W�i���u��&���9�2�������c �����GDM_qu�.9�FY3����c ���GDUgy/u�6/��UPDATES�.U ;/��FRS�:\S/�-o�Up�dates Li�st�/��PSRB?WLD.CM�/���"�/�/��PS_ROBOWEL�� g�\?n?���?���?�? W?�?{?O�?	OFO�? jO�?{O�O/O�OSO�O �O�O_�OB_T_�Ox_ _�_+_�_�_a_�_�_ o,o�_Po�_to�oo �o9o�o�ooo�o( �o!^�o��� G�k ���6�� Z�l�������C��� �y�����D�ӏh� ������-�Q���� �����@�ϟ9�v�� ��)���Я_������ *���N�ݯr������ 7�̿[�ſϑ�&ϵ� 7�\�뿀�Ϥ϶�E� ��i���ߟ�4���X� ��Qߎ�߲�A����� w���0�B���f��� ���+���O���s��� ���>���O�t��������$FILE_� PR� �����������MDONLY �1@���� 
 �5�Y�0}�= f/����O� s�>�bt �'�K��� /�:/L/�p/��/ �/5/�/Y/�/ ?�/$? �/H?�/U?~??�?1? �?�?g?�?�? O2O�? VO�?zO�OO�O?O�O�cO�O
_��VISB�CK������*.�VD_[_�@FR�:\F_�^�@V�ision VD file�_�O�_ �_�Oo�O)o�_:o_o �_�oo�o�oHo�olo �o�o7�o[m( � �D��z� �3�E��i����� .�ÏR��������� A�ЏR�w����*��� џ`����������O����MR_GRP �1A��L4�C�4  B�9�	 ��񝯯����*�u���RH�B ��2 ���� ��� ���ݥ���������ި�%�ߤA�5���_�J��KnI���HemT��b�R���P����M���q� F����HuEYG��:;��=;|���@W���@�ۡ�����E��� F@ %�5U1ŝ�J��N�Jk�H9��Hu��F!��/IP�s��?@�u��ÿ9�<9���896C'�6<,6\b����B���A���BZ��B����BkIA��u���#�HAx�ԫB3�nB6���A�SA��L��'ߚ�A9�A�?�M��r�ߖ߁���ߥ�  >����AE�5@5� �߯����4��X�C� h��y��������v��BH9� ��8�����҃�k��F��X�5�
��P�X�P�l�`�w������B�����M�@�3�3��������U�UU!U<�	>u?.�?!����k����=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7�:��7p��D�@ ?D�� C�@�U+C���Ώ�'�� �����-�/�C/� #/1��/Y�/�/�/�/ �/�/�/0??T???x? c?�?�?�?�?�?�?�? OO>O)ObOMO;�N� P�^O�OZO�O�O_�O +__(_a_L_�_p_�_ �_�_�_�_o�_'oo KoXi�Xo~o�o�oi� �o�o=o�o�oB T;xc���� �����>�)�b� M���q���������ˏ ���7�/{/%/7/ ��[/��/ܟ�� �� $��H�3�X�~�i��� ��Ư���կ���� D�/�h�S���w����� �O㿩�
ϥ�.��R� =�v�a�sϬϗ��ϻ� ������(�N�9�r� ]ߖ�]o�������߷o �{�$�J�5�n�U�� y������������ 4��D�j�U���y��� ������������0 T�-��Q��u��� ���ϟ5GP; t_������ �//:/%/^/I/�/ m//�/�/�/�/ ?ǿ !?�?Z?E?~?i?�? �?�?�?�?�?�? OO DO/OhOSO�OwO�O�O �O�O��
__._@_� d_�O�_s_�_�_�_�_ �_o�_o<o'o`oKo �ooo�o�o�o�o�o �o&J5nYk �k}����� 1��U����y��� ď���ӏ���0�� @�f�Q���u�����ҟ ������,��P�? q�;?��[���ί��� ݯ��:�%�^�I�[� �������ܿǿ �� �6��OZ�l�~�E_O� ������������2� �V�A�z�e�w߰ߛ� �߿�������,�R� =�v�a������� ���'�I�K��7� 9�?���o������� ����8#\G�k �������" F1jUg�g� �����/�/B/ -/f/Q/�/u/�/�/�/ �/�/?�/,??P?;? t?�?MϪ?�?�?���? Ok?(OOLO3O\O�O iO�O�O�O�O�O�O�O $__H_3_l_W_�_{_ �_�_�_�_�_o�_2o Do�eo/����oe��o ���o��
%o.R =vas���� ����(�N�9�r� ]���������ޏɏ� �׏8�ӏ\�G���k� ������ڟş���"� �F�1�C�|�g����� į�?ԯ�����?B� ��;�x�c�������ҿ �������>�)�b� M�_Ϙσϼϧ����� ����:�%�^�I߂� Io[o��o�ߣo�o� �o3��oZ�u�~�i�� ����������� �� D�/�h�S���w����� ������
��.��� �'�s���� ��*N9r ]������� /ۯ8/J/\/n/5��/ ��/�/�/�/�/?�/  ?F?1?j?U?�?y?�? �?�?�?�?O�?0OO TO?OxOcO�O�O�O�O����$FNO �����A�
F0Q� P T�1 D�|���@RM_CHKTYP  �@�����@��@��QOMP_MIN�"P����NP� � X�@SSB_�CFG B�E? ��{_���rS�_�_�ETP_�DEF_OW  ���-R�XIRC�OM!P�_�$GE�NOVRD_DO�CV���lTHR�CV dedd_E�NB�_ `RA�VC_GRP 19CdW�Q X�O�o �O�o�o�o�o�o& J1nUg�� �����"�	�F� X�?�|�c�������֏�������0�bRO�Up`I�HQP�����R��8�?T쀟3�|�����>��  Dڟl�l��@@�B�������o�4�g`SMT
mcJtm蕗�������AHOSTC]R19KO�pP�a�k M������0�  27.0zG�10�  e'� t���������b�ۿ�����4�˿ų	anonymous8� f�xϊϜϨ����л���%�'��[�0�B� T�f�x�ǿ�߮����� �Ϗ�E��,�>�P�b� ��������������� ��(�:���^�p��� �����������  $s�������� �����K� 2 DVh������� ��5GYkm7/ �v/�/�/�/�/�/ �/??*?M/��r? �?�?�?�	//-/O A?c/8OJO\OnO�O�/ �O�O�O�O�OOM?_? 4_F_X_j_�?_�?�? �__%O�_oo0oBo �Ofoxo�o�o�o�__ !_�o,>�_�_ �_��o��_��� �So(�:�L�^�p�� ��o��ʏ܏� �u�~١ENT 1LO�� P!��E�  A�3�p�_���W� ��{�ܟ���ß�6� ��Z��~�A���e�Ư �������� ��D�� h�+�=���a�¿��� ��
�Ϳ�@�/�d�'� ��KϬ�oϸϓ���� ��*���N��r�5ߖ� Y�k��ߏ��߳����QUICC0!����p�3�1q�M�_���3�2�����!ROUTER������`�!PCJ�OGa�<�!1�92.168.0�.10:��NAM�E !"�!R�OBOT���S_�CFG 1K"�� �Au�to-start{ed`tFTPkH���s��� ���$�'9 \J������ Jv!3E/Y{1/ b/t/�/�/g�/�/�/ �/?'/�/:?L?^?p? �?�?Qcu�?? O O/$O6OHOZO)?~O�O �O�O�O�?kO�O_ _ 2_D_V_�?�?�?�_�O �_O�_�_
oo�O�_ Rodovo�o�_�o?o�o �o�og_y_�_1 �o��_����� �o�&�8�J�mn�� ������ȏڏ);M _a�F��j�|����� ����֟����/�ɟ ßT�f�x�������� �!�#��W�,�>�P� b�t�C�������ο� ����(�:�L�^ϭ� ��ѯ������� � �$�6��Z�l�~ߐ� ����G�������� ����T_ERR �M��.�>�PDUS_IZ   �^����U�>n�WRD� ?��� � guest\��������������SCDMNGR�P 2NX����p��\��KM� 	P01�.14 8�� �  y��}�B�    ;����� ���߇�����������������~��\��������|���  �i  �  
����ҕ�����+��������
����l��.؋�"��luop �
dy�������&�_�GROU8�OM�� �	0�p�07��	QUPD  d��U��!TY��M�@�TTP_AUTH 1PM�� <!iPeOndan�������!KARE�L:*���K�C����VI�SION SET� ://���Q/?/ i/��/{/�/�/�/�/��/"?�/>YCTRL QM�P�v5���
��FFF9�E3.?��FRS�:DEFAULT��<FANUC� Web Server�:
Y��� A<OO*O<ONO`O<��WR_CONFI�G R<� ��?>�IDL_CP�U_PC�0��B�ȩ��@�BH�EM�IN�L���DGNR_IOG�|��S�@�NPT_SIM_�DOV[TPM�ODNTOLV >3]_PRTY)X�B��DOLNK 1SM����_�_�_�_�_��_o|RMASTE�P&|R_O_CFG"o4iUODEo6bCYCLEdo4d�0_ASG 1T<���
 o�o�o�o �o!3EWi{����k�bNUM�{�Q��08`IPC�H�o58`RTRY�_CN�0
RQ�6bSGCRN>{�Q�U�1 6ba`?bUM���p����$J23_�DSP_EN� �M�ᆀOBPROqC��LUMiJOG��1V�@Q�8G�?��{?Ń�POSRE��VKANJI_`d�
_HH��V�W�L}6h�<1�C�CL_L�@�r��H�EYLOGG+INB`���Q�P�LANGUAGE� �6�B�4 ,�>�LGW�Xf?��+����x% ���?���@���'0���`$�>MC:\�RSCH\00\��?�N_DISP YM�Ĩ�|�z��<�LOCGR�BDz��DA�OGBOOK Z�kR�P�T�X��B�T� f�x�����������v6	�<��⸥����_BUFF K1[�]� I�2�� H�S�h�d�n��ϒϿ� ����������+�"�4� a�X�j�|ߎ߻߲�����ߔ�ˀDCS }]� =��;� ��C��5Y�k�}����IO 1^�k t��� ������� ��� �2�D�X�h�z� ��������������
�0@Rdx��E^PTM  GdR2 ����0B Tfx����� ��//,/>/)Ĩ �SEV:����TYP���/�/�/ �-�RS�0��*�2��FL 1_��@��9�9?K?]?o?�?�?L�?�/TPѐ��"}ݭNGNAM���p�tU�UPS��G�I���E�A_L�OAD��G %���%��_MOV�[�aO�DMAXUALRM�w��x{@A�dQ:�<��C��y@C��`��Oj�lM�@̀�Ҁa�k �X�	V�!�p+e���O Τ,RX_C_U_�_7�|_ �_�_�_�_�_oo;o &o_oqoTo�o�o�o�o �o�o�o�o7I, mX�t���� ��!��E�0�i�L� ^�����Ï�����܏ ��A�$�6�w�b��� ����џ��������� �O�:�s�^������� ͯ���ԯ�'��K� 6�o���d�����ɿ�G�D_LDXDIS�A�0���MEMO�_AP�0E ?a+
 � ѹ%� 7�I�[�m�ϑϣ�y@�ISC 1ba+ �����'T,���
� ��C�.�g�Nߋߝ�� �߀�����	���?� ��N�"������ ��b������;�&�_� F��������x����� ��7��F �|���Z�� �3W>{���p���/��_MSTR ca-~%SCD 1d���m/��/|/�/�/ �/�/�/?�/3??W? B?{?f?�?�?�?�?�? �?�?OOAO,O>OwO bO�O�O�O�O�O�O�O __=_(_a_L_�_p_ �_�_�_�_�_o�_'o oKo6o[o�olo�o�o �o�o�o�o�oG 2kV�z��� ����1��U�@��y�/MKCFG �e--��<"LT�ARM_��f�;�� v���|���METPU��n���5)NDS?P_CMNT���8��#�&  g-.a��v���y���#�PO�SCF/�:�PR�PM.� �PSTOoL 1h��4@��<#�
��t���� �����/�q�S�e� ������ݯ��ѯ�����I�+�=��i�#�S�ING_CHK � ǟ$MODA�QӃi��a�����D�EV 	K*	�MC:�HSIZ�E�--ȹ�TAS�K %K*%$1�23456789� V�hŷ�TRIGw 1jK+ lK%3%�a���  ������M#8�YP#���5$���EM_INF� 1kڇ �`)AT&�FV0E0��a�)�I�E0V1&A�3&B1&D2&�S0&C1S0=>P�)ATZaߵ���H����p���	��A�9���]�D��� G߸�k�}ߏߡ�� ��6�m�Z�l���K� ����������� �� ����hs�-����� }����@R v);M_�� �+/*/�N/	/r/ �/k/�/[m�/�� �&?8?�\?�/�?;? E/�?q?�?�?�?O�/ 4O�/�/??�OA?�O �O�?�O�?_�O_B_�)_f_��ONITO�RJ�G ?��  � 	EXEC�1p��R2�X3�X4��X5�Xy��V7�X8
�X9p��R0Bd�R d�Rd�Rd�Rd�R d�Rd�Rdbdb�c2h2'h23h2�?h2Kh2Wh2ch2�oh2{h2�h3h3�'h3�R��R_GR?P_SV 1��>����(q���%I���SǾ!����h���(�>gr�+�@�_DR�&Λ�PL_NAM�E !��p��!Defaul�t Person�ality (f�rom FD) RR2-q 1m�)deX)dh��q7�X dv� �� $�6�H�Z�l�~����� ��Ə؏���� �2�D�V�h�t�2����� ��Ο�����(�:���<��d�v������� ��Я�����*�踝R,r 1r�yհ=\��, ������f� @D�  &z�?���f�?������A'�6z�ܿ���;�	l��	 ��xJ�԰�����˰ �< ���� ��IpK��K ��K=*��J���J���JV尻�"�ɱT���:�L�Ip@j��@T;fb��f��n���%�4��=�N����I���g��a������*��*  ´�  ��P�>��������n�?z����n���Jm���� 
�ғ�`%��Ī�9��� �`��  P}pQ�}p�}p|  ��r�/׈�+�	'� �� ��I� �  ��J��:�È��È=G�����6Ç�	����I  �n @
�+�l�$��l�!��9�A�7�N�p|�  '��_���@2��@���f�Z��@��C��C�p_C�@ C��C���C��o�
�A��q�   U@���
0ǉB�p*�A��2���0`�o�R�n�Dz��q���߁�������2���( �� -����������o�' ���!�o�M�� �?�ff ��/A�� ���v�7�a��
>N��  P��2�(o� �e�����ڳڴD�/?��o�x"Ip�<
6b<߈�;܍�<�ê�<� <�&�KNA둳��n�O�?fff?�?y&�3�@�.��J<?�`� M����.ɂ���� �lƴa2//V/A/ z/e/�/�/�/�/�/�/8�F�p�/4?�/�X?�y?�K?�?��E��� E��G+� F���?�?�?�O'OOKO6OoO.�BL��B�_0���O UO[��OcO_o?5_�?�\_�O�_�_�_�_U
��h��V�W>�r_on_/oo,oeoF�GA��d;���CRop�oNoD������o��o%5yķD��f8C|�spCH5�"Z�d����a�q@I��~N'�3A��A�AR1AO��^?�$�?���;��±
=���>����3�?W
=�#���{�e��n�@������{����<���~(�B��u��=B0�������	���H�F�G����G��H��U`E���C��+���I#�I���HD�F���E��RC��j=z�
I���@H�!H��( E<YD09ڏ�׏��� 4��X�C�|�g�y��� ��֟������	�B� T�?�x�c��������� �ϯ���>�)�b� M���q��������˿ ��(��L�7�Iς� mϦϑ��ϵ������ $��H�3�l�Wߐ�{� �ߟ߱��������2� �V�A�z��w��� ����������R�:�q(�q���������e��xv����a3�8���<���a4Mgs�������IB+���a?���{�&&	�fT�x���eP�P��A�O	\�`��*<��R^�p�����  ����*//N/</ r/�)�O� ��/�/�%�Q�/�/�/??'?9?  N?l/�?��?�?�?�?�2 wF�$�Gb��A��@a�`rqC���C@�oTO� q�{OF�� Dz@��� F�P D��aO�O�I�cO�O�O�__1_�c?��ͫ@@8Z^4� �� �� �n
 8_�_�_�_�_�_�_ oo+o=oOoaoso�o��zuQ ������1��$MSKCFMAP  R5� `6�uQqQ�n�cONREoL  ��a�� �bEXCFEN�Bw
�c�e qFN�C'tJOGOV�LIMwdprd��bKEYwsu��bRUNc|su��bSFSPDTY��p)vu�cSIGN|tT1MOTe�q�b_CE_G�RP 1sR5�c\:�I�2�m���D i���a�Ώ��Ï��� (�ߏ�^������K� ��o�ܟ��ɟ� H���l�~�e���Y�Ư�د�����F�`TCO�M_CFG 1tB�m�V8�J�\�
�__ARC_$r��2yUAP_CPL���6tNOCHEC�K ?�k �׸տ����� /�A�S�e�wωϛϭ��������kNO_WAIT_L�w�e��NT �u�kw[�5�_ERR!�2v�i�� ߠ߄�߾��c���ߴ�T�_MOc�wj�, ����3���PA�RAMd�x�k��tV#���=?�� �=@345678901��������� ���+�U�g�C�����y�������t����UM_RSPA�CE�olV>H�$?ODRDSP��v�2xOFFSET_�CART��yDI�S�yPEN_FILE� jq^�+�v��OPTION_I�O�YPWORK� y'�5s  x�fRuQ��2��2	 �	2���[ RG_DSBOL  R5sx\��zRIENTT5Op!C�oP�a�.A[ UT_SIM�_D��b�b[ V~_ LCT z?��*+^�)�_PEsXE�,&RAT8 �jv2u�p0"� UP S{.�PS0��/��/�/�/�)�$O�2� �m)deX)d�h��X d ��?-???Q?c?u?�? �?�?�?�?�?�?OO�)O;OMO_OqO�O�H2 
?�O�O�O�O�O__1_C_U_%�<�O_�_ �_�_�_�_�_�_o!o�3oEo�O� �Ov 1�r(���(���07�, ��lp�` @D��  �a?��c�a?m�a%�D�c�a����l;�	l�b	 ��x�J�`�o�u��` �< �	p�� �r��H(���H3k7HSM�5G�22G���Gp
������c�Yk|��CR�	>��qȋs�a�����*  ���4�p�p��pT����B_����=j%��t�q� )�/��aD�����~�6  ���UP� Q� �� |�Б�������	'�� � ͂I�� �  ��i�=���������a	���I  �n @)��m�C���m��[��N���  '� ��~q:�pC�C�@�s�p�C���ҟ 5�
���=x@#�7~H9�^�n�B�I�A��Q��� 0�q��bz比������ȯ�����( �� -݂*�΁6���Am� �0rx���m�lp �?�fAfU ܫN�`�����n�8m྿̺>N�  P�aզ(m� ������ q�c�d#/?��m�xA�n��<
6b<߈�;܍�<�ê�<� <�&1j�m�A0��c��ƾn�?fff?0�?y&����@�.���J<?�`�� l�����dѩ�e�ϟg ߋ��d��Q�<�u�`� �߄߽ߨ�������� )� �M�8�q���
���j���f�E�� E��0�G+� F� ������ �F�1�j��U���y�[bB��A ��|����t�z��� 3��T��{����x��t��h��u�w�>��*�`N9K���A��Z�_�Cq�mc��?��//D///
T)���pٞ�a�`#CHT/A
$� !��!@Iܝ�'��3A�A�AR�1AO�^?�$��?�����±�
=ç>�����3�W
=�#��>��+e�� �������{�����<��.(��B�u��=�B0�������	3�\*H�F��G���G���H�U`E����C�+�Y-I#��I��HD��F��E���RC�j=�>
�I��@H��!H�( E<YD0X/�?O�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_s_^_�_�_�_�_ �_�_o�_ o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV h������� �1�C�.�g�R���v� ����ӏ��Џ	��-� �Q�<�u�`������� ϟ���ޟ��;�&��8�q�\�(�����,�����]��������p!3�8����ӯp!4Mgs8����IB+�+���a���{� E�E���s�����Ϳ��J�Pe�P���(�{�4��I�[�իR}Ϗ��ϳ�������  ���˿I�7� m�[ߑ��H� �������������p"�4�F�X�  mߵ���������2� F�$�Gb	��ϲ����!C���@�s�����~ F� Dz/���� F�P DC�����������,>P�?̯��@@W
}�R���������
 W���� &8J\n�p���*� �������1��$PA�RAM_MENU� ?q���  DEFPULSE��	WAITTM�OUT+RCV�/ SHEL�L_WRK.$CUR_STYL ;G,OPT]�]/�PTBr/l"CB/R?_DECSN � �,�/�/�/
???)? R?M?_?q?�?�?�?�?��?�USE_PR_OG %�%�?\#O�3CCR ���6G_HOST !�!;DxO0JAT�BO�C[OmA�C|�O/K_TIME"ܜB�  �GD�EBUG�@��3G�INP_FLMS�K�O(YT��9_*UP+GAUP \��g[�CH6_'XTYPE
����?�?�_o o#o5o^oYoko}o�o �o�o�o�o�o�o6 1CU~y��� ����	��-�V��Q�c�u���*UWOR�D ?	{]	�RS��	PNS2W�V$ڂJO�!���TE�@�VTRA�CECTL 1|vq�� ��_� ����|4��DT Q}q��c�(�D � _ L� p�QMt�� v�O� �o��� � ��� ������p��� p�Òp���w��Pv�� �v�� v�t�t�	�t�
t�t�t��t�t�t��@v��t�t�t�t�(t�V�v�t�t����v�t���v�� v��t�t��v�N�v�!�t�"t�#t�'�v�%�t�&t�'t�(t�)�t�*t�@�v�,t�-�t�.t�/t�0t�1�t�2t�3t�4t�5�t�6t�7t�8t�9�t�:t�;t�<t�=
t�>t�?t�n v�]� v�� v�� v�Dt�Z �v�Ft�Pv�Ht�It�Jt��Pv�s���7��@6�Q4Ĥ�6��6�T 6�U4�V4�W4�UX4�Y4�Z4�[4�U\4�]4�^4�_4�U`4�a4�b4�c4�Ud4�e4�f4�g4�Uh4�i4�j4�k4�Ul4�m4�n4�o4�Up4�q4�r4�s4�Ut4�u4�v4�w4�Ex4�y4Ĳ�6�{4� ����������ב�� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�l�Е ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ Е���_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
���_@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/�:/L/^/h!�$PG�TRACELEN�  g!  �_�f �|&�_UP ~�����!� �!�� |!_CFG ��%�#f!�!���$� �/�/;�"DEFSPD ��,�1�� �| IN~� TRL ��-�f 8�%G1PE__CONFI� ��%���!�$�<LID�#��-~�4GRP 1��7�!�g!A ����&fff!A+�33D�� D]�� CÀ A@6B1�f d�$I&I��1�0� 	 p?�"�+@O ´yC[ODKB|@�A�OmOO�O�O�Of!>�T?�
5�O4_F^0_� =��=#�
K_�_G_�_�_�_�_ �_c_�_&o�_6o\oGo�  Dz�c�of 
 qo�oao�o�o�o�o 0T?xcu������IK
V�7.10beta�1�$  A��E/�ӻ�Ay f ,�?!G�C�/>��+���0T����+�BQ�c�A\i�T�D;�{�p�"�B������Ə؏�T�O'O�2�8��\�G���k� ������ڟş���"� �F�1�V�|�g����� į���ӯ���	�B� -�f��ov���K����� �������>�)�b� M�rϘσϼϧ�����<�=�F@ �� '�۫%Wك�W߉ߛ� �6���������%� �I�4�m�X��|�� ����������3�� W�B�{���x������� ������S~� w�8����� �+O:s^ ������
�<�/ /R�d�v�l/~/�ߥ/ ��������/�#?5?  ?Y?D?}?h?�?�?�? �?�?�?�?O
OCO.O gORO�O�O�O�O�O�O �O	_�O-_?_jc_u_ $_�_�_�_�_�_�_�_ oo;o&o_oJo�ono �o�o��(/�ob/ P/&Xj�/��/�/ �/�/��o��3�E� 0�i�T���x�����Տ ��ҏ���/��S�>� w�b�������џ���� ���+�V_O�a���� p�����ͯ���ܯ� '��K�6�o�Z����o �o�o޿*<n D�rk�}Ϩ��� �φ������
�C�U� @�y�dߝ߈��߬��� ������?�*�c�N� ��r��������� 0���;���_�q�\��� �������������� 7"[F����ο ����(�0^� Wi�Ϧϸ�v�r ��/�///S/e/ P/�/t/�/�/�/�/�/ �/�/+??O?:?s?^? �?�?�?�?�?�?�O 'O�?KO6OoO�OlO�O �O�O�O�O�O_�O_ G_2_k_����_�_ �
ooJCoUo ����oL_�o�o�o �o�o?*cu `������� ��;�&�_�J���n� ����ˏݏO�� 7�"�[�F����|��� ��ٟğ���!��� W��_�_�_�����_�_� o���6b�$PL�ID_KNOW_�M  bd��j�#�SV ��3e=�:e��z�����7��¿������j�vmC�M_GRP 1�P���`d�bd@I�߶B�_�
�_��� ��t��@ǘϾ�^��� �ϮϪ�
�����F�� d�(�Zߠ�^����ߔ� �����*��� �f�$� L��Z�|���������,�>�#�MR'Éb.�Tg��� � ���������������� ����Q+%7�� �������� M'!3��������Y�ST'�1W 1�3e3 �i�;0:o A >/g� </N/`/r/�/�/�/�/ �/�/�/?C?&?8?y? \?n?�?�?�?�?�?	O�'2(.:/j��	<=O.3'O9OKO]O�!#4vO�O�O�O!#5 �O�O�O�O!#6_&_8_J_!#7c_u_�_�_�!#8�_�_�_�_!#M_AD  wd3#�x`$PARNUM  ++�5o"WSCHOj ]e
�gppa�i=��eUPDpo��e�t"_CM�P_$�R`ؠ`'�;�)tER_CHK7u��;�Or4F{�RS|�2�#�_MO�Q`��u_�be_R/ES_G' �+-O ���H�;�l�_��� ����Ə���ݏ����w&@�|�5��u u@R�q�v��s�@���� ���sPП����sbP �.�3��s�PN�m�r���s `�������rV �1�P���b@cX���p�$@cW��(��(�@@cV��4���rTHR_�INR|�Taud�<�MASSI� Z�]�MNH�{�MON�_QUEUE Q�.�bvg��g�bdN.pUrqN��`{ΰ�ENDб��EX1E����`BE��ڿ>˳OPTIO׷�{�ΰPROGRAM7 %��%Ͱ���o̲TASK_I�Qd@�OCFG Ꭾ��o����DATuAe���@�2�N�`�r߄ߒ�<� �������ߖ��!�3�xE�W�
�INFOe��"ݘ������� ������)�;�M�_� q����������������n�z�"� �!���OpDIT ���s�WERF�L��#RGADoJ �b
A��0��?��P��IOORITY��av��MPDSPX��eU����OG$ �_TG� K���ET�OE��1�b _(!AFD�E�p���!tcp|��!ud�>�?!icm��nFXY_���b{���)� *J/\/` ���G/�/k% w/�/�/�/�/�/?�/ 2??V?h?O?�?s?�?z�?*�PORT3��Rc���u�_CARTREP�|bk@SKSTA��^�zSSAV���b
�	2500H8�63(�ς5D1�*b`@�����s�O�O�G	PURGE��B�	�yWF�@DO��$�evW�T�a��:WRUP_DE?LAY �bT�R_HOT{��%�o�_TR_NOR�MAL{�}_�_�VS�EMI�_�_oCaQ�SKIP1��u�Cx 	bO\o\@ Jo�o�o�ojh�u�o�g �o�o	�o?-O u��_���� ���;�)�_�q��� I�������ݏ��Ǐ %��I�[�m�3�}������ǟٟ�ͥ�$R�BTIFR�RCgVTM.+D�	��DCR1c�8l����C�CB���C�7?����=>�<�Wem��=��x\A��yv�?�jݼ��1ho���dn<
6b<�߈;܍�>u�.�?!<�&ǯ���)�ŰH B�T�f�x��������� ҿ������>�)� b�Mφ�qσϼϟ��� ��5��(�:�L�^�p� �ߔߦ߸��������� ���6�!�Z�E�~�� s����	������ � 2�D�V�h�z������� ��������
��. RdG����� ��*<N` r�o����� /�&/	//\/��/ �/�/�/�/�/�/�/? "?4?F?X?C/|?g?�? �?�?�?�?�?�?O0O s/TOfOxO�O�O�O�O �O�O�O__,_OP_ ;_t___�_�_�_�_�_ �_oGO(o:oLo^opo �o�o�o�o�o�o�o�_ �_$H3lW� ����o�� � 2�D�V�h�z��������ΈB�GN_AT�C 1�O� �AT&FV0�E0΋ATD�P/6/9/2/�9�ATAΎ�,AT%G1�%B960�W+++3�,.�Hc��,B�IO_TYPOE  �����ЏREFPOS1� 1��� x	��������?� P����6�������V��߯z���� �9�Ǜ2 1�����$�ࢿ �ƿD�ё3 1�^�p�����:�%�^�>ܿS4 1�����Q��Ϻ���q�S5 1��ϚϬ���d��O߈��S6 1� �/�A�{�������S7 1����������y��0�S8 1�G�Y�k��#���G���SMASK ;1���  
����Ne�XNO��;�A������͑MOTE � ��ʔ��_CFG� ���<���̒P?L_RANG���q���POWER ��^ ��SM_�DRYPRG �%��%��dTA�RT �V�
U?ME_PROs�� ʔ_EXEC_?ENB  =���GSPD� #���4TDB>PRM\_PMT_m�TQ �����OBOT_NAME ����׉OB_OR�D_NUM ?�V��H8�63  �t /��!\<� { # 	r*!7@�"D|<����PC_TIMEO�UT6 x��S2�32
1�� �LTEACH PENDAN_ ����e�����Maintena�nce Cons��r���*"�/�KOCL/C� :����/? No Usee��/U?��v#NPO218�����t!CH_�L� ���7�	��1�;MAVAIL��a#�������SPACE1 2�ٜ �?%dH�9��eF%�<��L8�?H �9�O�?�O �O_�O(_#WTOfOxO �O8_�O�O�_�_�__ o i��4mT_f_x_ �_�_�_�_�o�o�oo� .�5;A2@N ROdovo�o6�o�o�����4��I�N{3 ]o���S��� ���ޏ0�Q�8�f�N{4z�������p�� ��8���M�n�U���N{5������͟ߟ�� �%�4�U��j���r���N{6��Ưد��� �� �B�Q�r�5χϨ��Ͻ�N{7ѿ���� ���=�_�nߏ�Rߤ��߬���N{8�� �� $�6���Z�|ߋ��o����������N{G ���� ���$
�� C�e#p��� ����������:hL���@2��+��^�!dt  Y�k������� ��8oR~ q������/ /=/7Ikm�/ ���/�/�/??+?�=?3/]?W/i/�/�=; `�� @NP�5@<�?�/�) A�5�? 1OCOI?#J$OVO�O�O �O~O�O�O_�O�O�O _^_ _2_D_v_�_�_ �_�_�_o$o�_�_
o<o~o@oN<
O�oN{�_MODE  �+��iS �+��ox?v:_��?'y�z	��o�CWO�RK_AD�m�{_�q�R  +������p_INOTVAL�`@�z�R_OPTION�1� u��VA�T_GRP 2��+�]�(���L��ԏ� ��
��.�@���d�v� ��O�o���dX�ß� ���ϟ1�C�U�g�)� ��������ӯ�{�	� �-���c�u���I� ����Ͽ��ϛ�� ;�M�_�!σϕϧϹ� {�������%�7��� [�m��Aߏߵ����� �����!�3�E�W��� {����s������� ����/�A�S�e�w��� ����������� +��Oas��� ?����'9�K[����e��$SCAN_TI�M�a��\��R ��(�30(��L8z�J�p�p
WtZ��2#Nq!�#Y�:.(/V1�#M"2{$D!!d�(~!�!�r #])�0��/�/�/��r�)�/  P5u�0�2  8��?U?g?>1D�� j?�?�?�?�?�?�?�?�O#O5OGO?Nq�%�RO�O�O[N![q;�o�t�Nq�p]M�t���Di�t!c{  � lM"Nq�A!
%� 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�gS �o�o�o'9K ]o������ ���#�5�G�Y��o �o�K������Џ�� ��*�<�N�`�r��� ������̟ޟ����1�  0�B|�_ g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ�p�� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑ��� ����������0�B� T�f�x�������� ������,�>�P�J�V�  �1�������� ��������1C Ugy�����8��	 �y3 "HZl~��� ����C&5/�</+&�r! �5/q-	1234�5678R�+��L{0�@�/ �/�/�/�/?3,? >?P?b?t?�?�?�?�? �?�?'OO(O:OLO ^OpO�O�O�O�O�O�? �O __$_6_H_Z_l_ ~_�_�_�_�O�_�_�_ o o2oDoVohozo�o �_�o�o�o�o�o
 .@Rdv�o�� ������*�<� N�`����������̏ ޏ����&�8�g�\� n���������ȟڟ����"�+&s�C�U��:�Z��������C�z  Bp  � ���2/$@���$SCR_GRP� 1�(�e@(�l�� �@ Z! �U!m�	 #�-�=� 6�n�p�l�S�y(J�w��e������3%D!ʰ֠o��ป���M-10i�A 890�%90�� Ɓ M61CA �#�-I���#�
\�l�,�O'|�Z!�S�;�o�}�	n������������X � ,���Y"N�a����ߖ� i�@�.!`/��m�����\"��B�Š�J��H�a�H�A֠p�  !@. ��l��?����D�HŠ���H�F@ F�`����� ��;�&�K�q�\��� ����<�����������B���YD }h������ �
CҾ?4#��0/v/�%��
��������V�j�@����/ B�*'���P���EL_�DEFAULT � C�����X!MIPO�WERFL  �P�p%W"} WFDO�e& p%��ERV�ENT 1����I�n#=�L!DUM_EIP���(�j!AF_�INEd ?�!�FT�/7>�/[?!�K߀? �J?�?!�RPC_MAI�N�?�8��?�?�3V�IS�?�9��??O!7TP2@PU6O�)�d.O�O!
PMON_PROXY�O��&ezO�ORB�O�-f��O#_!RDM_�SR��*g_o_!#RL(�_�$h^_�_K!
�0M�O�,i�_�o!RLSYN�Co.i8�_So!�ROS�/zl�4 Bo�on?�o2S�o�o�o �o5�oY }D �hz����� 1�C�
�g�.���R�����'ICE_KL �?%�+ (%SVCPRG1�� ������3$�)�"�4L�Q��5t�y�"�6�����7ğɟ��=��/�9�� 脆_A���i��� ���>����f��� ��	�끶�1��ޟY� �����.����W� ѿ�������!�� ϯI����q����� �G����o������ ����9�;�翹�˂ �ҏ䀄���á���� ��� �9�$�]�H�� ��~����������� #��5�Y�D�}�h��� ������������
 C.gR�v�� ���	�-Q cN�r�������/)//M/��_�DEV �)��MC:U(���]g$OUTYB�`!x&c(REC 1q���` �  ` _ 	 ` ` ` ` �!�!U+�#���U/�.�$1��"?`!` 8�:
 �P�b�6 s�'� � �  '� _�  =0f�ը�"�#�!� ` /J` �` ��=y �y }�y �����` B� D�?O�%��|0���<S  ��iH� �0_��?� O�` �4)�` ��?��`!y �*�0�` k� NPO�OVOc݀;[0�0~�1o  �� �i�O !� � �j04,` �xO��y )��!�Dn� M�O]_��Oc��O�@�F� �O
__._@_R_d_I�f�6r _�H�i@�4�x�C�@�,�_�!r` �` C`m �P#�_�fy U�y �y �y �<1�To�ooh$0k ��  � �1  W �i@=�o ;@غ2�0�   K`$V|o�dy �y �y �Dq��! a�oh[��l�0k`�bR  �Ȣ lP
5�2j` �` �(�c�4���D��!��t~�kj�0k� ��3���`  #"T�j2;� ` L` ��� wO���y �y ��qy ��QX����taĀ<Đ?g ���?�?�?�?��ď"F� �;T�f�4����'�+�` =� �T� ��
` Q� ,�������H��` U� F���x�02y0 �  �T�B�x�f������� ү������,��P� >�t���h�����ο�� ޿��(�
�8�^�L� ��pϦϔ����Ͼ� � ��$��4�Z�H�~�`� rߴߢ��������� � 2��V�D�f�h�z�� ��������
���.�� R�@�b���j������� ������*<` N�r�����%oV 1��, P 8�� :���*X  p� 
t�pJc(�TYPE�/e"HE?LL_CFG���&�� ��"�� %RSH��// </'/`/K/�/o/�/�/ �/�/�/?�/&?8>�pr:>����` %K?@y?�?F=J1J1�p gA��=�1�p��a22�!�d�?�?�HK 1���a�?AO<O NO`O�O�O�O�O�O�O �O�O__&_8_a_\_�n_�_|OMM ��_FTOV�_ENO�nwO�W_REG_UI��__IMWAITp�Rq�6kOUTf� iTIMe��ZoVAw�1o#a_UNIT�S�fw�MON_ALIA�S ?e�Y ( he�o�o 0��o]o��> ������#�5� G�Y�k��������ŏ ׏������1�܏B� g�y�����H���ӟ� ��	���-�?�Q�c�u�  �������ϯᯌ�� �)�;��_�q����� ��R�˿ݿ��Ͼ� 7�I�[�m��*ϣϵ� ���τ����!�3�E� ��i�{ߍߟ߱�\��� ��������A�S�e� w��4�������� ��+�=�O���s��� ������f����� '��K]o�,� �����#5 GY}���� p��//1/�U/ g/y/�/6/�/�/�/�/ �/�/?-???Q?c?? �?�?�?�?�?z?�?O O)O�?:O_OqO�O�O @O�O�O�O�O_�O%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3o�_ Woio{o�o�oJo�o�o��o�o�c�$SM�ON_DEFPR�O ����4q �*SYSTEM*� . "vREC�ALL ?}4y� ( �}5xc�opy fr:\�*.* virt�:\tmpbac�k}q=>desk�top-b25t�4o0:5440� �r����z}6tua|��w�<�N���:uts:ord�erfil.da�t�����͏ߏ}=1urmdb:��� &���8�J�\��qs� ����̟ޟ����� '�8�J�\�o���
��� ��ȯگ�����#�4� F�X�k��������Ŀ ֿ������0�B�T� g�y��Ϯ������ �������>�P�c�u� ϙ�+߼���a������)�:�L�^� }
�xyzrate 61 ���#���������!t��15432 ���9�K�]���1���!����������7��:prog�ram_1.tp��empߏ���= Ob�����*�� �r�� �9K] ���&���n ��5/G/Y/�� /"/�/�/�/j|� �/1?C?U?h/��/?�?�?�?��;tφ�~? �3/OAOSO��2��O �<'O�O�O�O���ߏ� �8�O<_N_�O7��_ _�0-_�_�_�?�?O �_+_<oNo�_sOo�O )o�o�o�o�O�_�o'_ 8J\o_ �_� ��m���4�F��X�k?}?:16056�?'���ʏ܏o/�� ����6�H�Z��/�/? �,���ϟ�t��� ��;�M�_��_o�o� ����ӯfoxo������8�J�\�j��$SN�PX_ASG 1߼������ P 0 �'%R[1�]@1.1`���?�j�%��ֿ����ݿ �0��:�f�Iϊ�m� ��ϣ���������� �P�3�Z߆�iߪߍ� �����������:�� /�p�S�z������ �� ���
�6��Z�=� O���s����������� �� *V9z] o�����
� �@#JvY�} ����/�*// /`/C/j/�/y/�/�/ �/�/�/�/&?	?J?-? ??�?c?�?�?�?�?�? �?O�?OFO)OjOMO _O�O�O�O�O�O�O�O �O0__:_f_I_�_m_ _�_�_�_�_�_o�_ oPo3oZo�oio�o�o �o�o�o�o�o: /pSz���� � ��
�6��Z�=� O���s���Ə���͏ ߏ ��*�V�9�z�]� o��������ɟ
�ퟀ��@�#�J�v�Y�r�PARAM ����� �	��z�P��j�O�FT_KB_CF�G  ����ѤP�IN_SIM  �Ʀ�)�;�ɠ�r�RVQSTP_DSB �Ƣw������SR ���� & �������ΦTOP_ON_�ERR  �����PTN z��Aݲ�RING_PRM�� ��VDT_?GRP 1����  	ʧ��\�n� �ϒϤ϶��������� %�"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�w�t����������� ����=:L^ p������  $6HZl~ �������/  /2/D/V/h/�/�/�/ �/�/�/�/�/
??.? U?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFomojo|o�o �o�o�o�o�o�o3�0ѣVPRG_CoOUNT�����^rENB)�YuM��s㤐_UPD �1��8  
 G�����'�"�4� F�o�j�|�������ď ֏������G�B�T� f���������ןҟ� ����,�>�g�b�t� ��������ί���� �?�:�L�^������� ��Ͽʿܿ���$� 6�_�Z�l�~ϧϢϴ��������VuYSDE�BUGhp�p���d��y�SP_PAS�ShuB?.�LOoG ��u�s������  ���q��
MC:\xZ�
�[�_MPC`ݐ�u�����q��� ��q��SAV �bc��ԛ������SV�TEM_T�IME 1��{+ (�p֪t���s��N|T1SVGUNYS�piu'�u����ASK_OPTICONhp�u�q�q���BCCFG Ō�{I� B��5�`5�;zC�l�W�i� �������������� 2D/hS�w� ����
�.�R=va���� ����/��B/ -/f/Q/�/�/��  �/�/�/�/�/ ??D? 2?T?V?h?�?�?�?�? �?�?
O�?O@O.OdO RO�OvO�O�O�O�O�O _�H�_,_J_\_n_ �O�_�_�_�_�_�_�_ o�_4o"oXoFo|ojo �o�o�o�o�o�o�o B0Rxf�� �������>� ,�b�_z�������Ώ L�����(��L�^� p�>���������ܟʟ �� �6�$�Z�H�~� l�������دƯ���  ��D�2�T�V�h��� ��¿x�ڿ�
��.� ��R�@�bψ�vϬϾ� �Ϟ�������<�*� L�N�`ߖ߄ߺߨ��� ������8�&�\�J� ��n��������� ��"�ؿ:�L�j�|��� ����������� 0��TBxf�� �����> ,bPr���� ��/�//(/^/ L/�/8��/�/�/�/�/ l/? ?"?H?6?l?~? �?^?�?�?�?�?�?�? OO OVODOzOhO�O �O�O�O�O�O�O_
_ @_._d_R_t_v_�_�_ �_�_�/�_o*o<oNo �_ro`o�o�o�o�o�o �o�o8&\J ln������ �"��2�X�F�|�j� ����ď��ԏ֏�� �B��_Z�l������� ,�ҟ������,���J��$TBCSG_GRP 2����  ��J� 
 ?�  u���q�����ϯ ��˯��)�;�N�U���\�d, ��j�?J�	 HC�=�8�>����9�?CL  B�m���ܰ�z��β\})��Y  A�f��B�;��Bl��=�,�ɐ�Z�,��  D	�{�F�`�j�ACs��όϦϰ̖���@J��+�>�Q�� .�|ߙ�d�v���������؈J�	V3�.00m�	m6;1c��	*,�$�I�;�D�>���J�(���� r�D�s� ; #����D�����N�JCFG -��f� i�������������7�E��E�k� V���z����������� ����1U@yd ������� ?*cN`�� ����m����/ "/�U/@/e/�/v/�/ �/�/�/�/	??-?�/ Q?<?u?`?�?�?J�6� �?��?�?�?*OONO <OrO`O�O�O�O�O�O �O�O__8_&_H_J_ \_�_�_�_�_�_�_�_ �_o4o"oXoFo|o�o ���o�obo�o�o�o B0fTv�� �~�����>� P�b�t�.��������� ̏Ώ����:�(�^� L���p�������ܟʟ  ��$��4�6�H�~� l�����Ư���د��  ��o8�J�\����z� �������Կ
���.� @�R�d�"ψ�vϬϚ� ����������<�*� `�N߄�rߨߖ߸ߺ� �����&��J�8�n� \�~���������� ��� �"�4�j�X��� |�����n��������� 0TBxf�� �����, P>t���d� ���/(//L/:/ p/^/�/�/�/�/�/�/ �/? ?6?$?Z?H?j? �?~?�?�?�?�?�?�? OO OVO��nO�O�O <O�O�O�O�O�O_
_ @_._d_v_�_�_X_�_ �_�_�_�_o*o<o�_ oro`o�o�o�o�o�o �o�o8&\J �n������ �"��F�4�V�|�j� ����ď������O� $��O��f�T���x��� �����ҟ��,�� ��b�P���t�����ί ௚�����(�^� L���p�����ʿ��ڿ  ��$��H�6�l�Z� |�~ϐ��ϴ������ ��2� �B�h�Vߌ�� 8�����rߠ�����.� �R�@�v�d���� ����������N� `�r���>��������� ���� J8n \������� �4"XFhj |������/ 0/��H/Z/l//�/�/ �/�/�/�/�/??>? P?b?t?2?�?�?�?�?��?�>  @
C� 
FO
B�$T�BJOP_GRP� 2��5�  ?�
G�6B=C�DL��0��xJ�@�
D@ �<� ��@�
D� @@UB	 ��C�� �Fb  �C�VGUAUA>��1��E�E�I>��@�A��33=�C�L�@fff?�@?�ffB�@Q�E-_�8W�N��O>��nR\)�O�@�U����;��hCY��@�  @�@UAB�  A�$_�_�S~�UC�  D�A8�LwP�RO�z_�S�b��
:���Bl�P��P�D�Q�_�So
AAə�A��hcZQDXg�F�=qq�e
o�@�p��b��Q�;�A}Ȱ@ٙ�@L�CD	x`�`�o�ojo|o>B�\u�oh�Q�ts�a@33@QV@C��@�`exw�o>��D�u�*�@� p�qP<{�Nr�@@�PZv_p ����&�:�$�2� `���l�&���ʏ�� ��!�����@�Z�D�R�(����DT�
Fґ�E	V3.00�C�m61c�D*����DA
�� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I�&�CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;'`;Q���8�`F�O���
F��Q��K�2D�ESTPARS c �8O@3CHRe�ABLE 1�DKI.�
CP�%� ~ �P�P�P�	GA*P�	P�
P�P����
AP�P�P�N|�RDI��NA��@��¿Կ���`�Ohπz˄ϖϨϺ��΀�Sf�LC *ʍߟ߱��� ��������/�A�S� e�w��������� )Me�iߘ�$���1� C����%�7�IȀ�~
�NUM  �5�NA�@@ ���[���_CFG ������A@6@IMEBF_TTk�p��LCx�5VERY��6�K5R 1ОDK
 8�
Bd@� �0/�  � ������  2DVhz��� ��/�
/S/./@/�V/d/v/u_��b@�L
6@MI_CH�ANA L �#DOBGLVPCL�5A� ETHERA�D ?�550��M��/�/N?0F� R�OUT_ !DJ!��4�?q<SNMA�SK*8LC;125�5.�5��?�?2DO�OLOFS_DI�k��%9ORQC?TRL �mK���hM8WO�O�O�O�O �O�O�O
__._@_��|ON_`_�_a�PE_�DETAI8-JP�ON_SVOFF�#O�SP_MON ��J�2�YST�RTCHK ��DNg?�RVTCOMPAT�X53�T�P�FPROG %�DJ%	qaRAM_�17o�\APLAY�l��Z_INST_�M�0 �l�W�dUqS_WoibLCK�l��kQUICKMEx� #ibSCRE@p�-:tps��ib�a[p`y�"qp_�uy��Ti9SR_G�RP 1�DI ؕ�0��z����5�#�Y�G�� 2 ����S��o����܏ ǅ����)��M�;� q�_�������˟��ݟ��7�%�G�m�	�1234567�堃���b�XZu1���{
 �}ip�nl/ՠgen.htm�����*��<�R�Panel setup@�}6o��������ȿڿ o�e��$�6�H� Z�l�㿐�ϴ����� ����߅ϗ�D�V�h� zߌߞ��C�9����� 
��.�@��d��߈� ��������Y�k�� *�<�N�`�r����� ����������8 ��\n����-��nUALRM�`G� ?DK
   �	L?pc �������/�/6/�SEV  ��h&�ECFG ��]�&��}A�!   Bȣd
 7/�c-5�/�/ �/??%?7?I?[?m?�?�7t!�r��[ P�3ȏ�?B'Imf?wk�P(%*/O`
OCO .OgORO�OvO�O�O�O��O�O	_�O-_�<�d ��=�?;_I_?pH�IST 1��Y � (�  ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,�o�_�_oo �s� �_�]936�_ lo~o�o�o1b�o�o�o �o%�oI[m ��2���� �!��E�W�i�{��� ����@�Տ����� /���S�e�w����������L��QL����� �1�C�F�g�y����� ����P����	��-� ?�ί�u��������� Ͽ^����)�;�M� ܿqσϕϧϹ���Z� l���%�7�I�[��� ߑߣߵ�����ğ֟ �!�3�E�W�i�lߍ� ���������v��� /�A�S�e�w������ ����������+= Oas���� ���'9K] o������ �����5/G/Y/k/}/ �/��/�/�/�/�/? �/1?C?U?g?y?�?�? ,?�?�?�?�?	OO�? ?OQOcOuO�O�O(O�O �O�O�O__)_�OM_ __q_�_�_�_6_�_�_ �_oo%o/"/[omo o�o�o�o�_�o�o�o !3�o�oi{� ���R���� /�A��e�w������� ��N�`�����+�=� O�ޏs���������͟ \����'�9�K�6o���$UI_PA�NEDATA 1��������  	�}�]�����ȯگ��� ) �$�ᔒ�O�a�s� �������Ϳ���� �'��K�2�oρ�hπ�ό����������� Ha$�7�<�N� `�r߄ߖ��Ϻ�-��� ����&�8�J��n� U��y��������� �"�	�F�-�j�|�c�������������� +=��a�߅ �����F �9 ]oV�z �����/�5/ G/����}/�/�/�/�/ �/*/�/n?1?C?U? g?y?�?�/�?�?�?�? �?	O�?-OOQOcOJO �OnO�O�O�O�OT/f/ _)_;_M___q_�O�_ �_?�_�_�_oo%o �_Io0omoofo�o�o �o�o�o�o�o!3 W>{�O _�_�� ����pA��_e� w���������&���� ܏� �=�O�6�s�Z� ��~���͟���؟� '���]�o������� ��
�ۯN����#�5� G�Y�k�ү��v����� ׿�п���1�C�*� g�Nϋϝτ���4�F� ��	��-�?�Qߤ�u� �����߽�������� l�)��M�_�F��j� ������������`7��[�����}�l�@������������)�� $��Pbt�� ������( L3p�i������ /(������$UI_PANELINK 1����  ��  ��}1�234567890Y/k/}/�/�/�/�$ ��W/�/�/??+?=? �/a?s?�?�?�?�?S9�S *�=��U   �?O(O:OLO^O�? \1O�O�O�O�O�O�O �O_(_:_L_^_p__ ~_�_�_�_�_�_�_�_ $o6oHoZolo~oo�o �o�o�o�o�o�o
2 DVhz$��`���
�E0,/ A�M�/�p�S������� ʏ܏�� ��$�6�� Z�l�O����<�?���� �T!���1�C�U� g�Z3��������ǯٯ �z��!�3�E�W�i� �<��������C��ÿ տ����Ϥs5�G� Y�k�}Ϗϡ�0����� �����߮�C�U�g� yߋߝ�,��������� 	��-��Q�c�u�� ���:��������� )���M�_�q������� ��(�����~���7 I,mb��� ����3ƞ�� ��՟w������� �/��,/>/P/b/t/ �//�/�/�/�/�/? ?������^?p?�?�? �?�??��?�? OO$O 6OHO�?lO~O�O�O�O �OUO�O�O_ _2_D_ �Oh_z_�_�_�_�_�_ c_�_
oo.o@oRo�_ vo�o�o�o�o�o_o�o *<N`��� ������� �8�J�-�n���c��� ��ȏڏI��m"�� F�X�j�|��������/ ֟�����0���T� f�x�������?/?A? �o��,�>�P�b��o ��������ο�o�� �(�:�L�^�p����� �ϸ�������}��$� 6�H�Z�l��ϐߢߴ� �������ߋ� �2�D� V�h�z�	������� ����g�.���R�d� G���k����������� ����<N1r� ���;�� &8J=�n��� ���i�/"/4/ F/X/ǯٯ믠/�/�/ �/�/�/?�/0?B?T? f?x?�??�?�?�?�? �?O�?,O>OPObOtO �O�O'O�O�O�O�O_ _�O:_L_^_p_�_�_ #_�_�_�_�_ oo$o �_HoZolo~o�o�o� �o�og�o�o 2 VhK�o��� �����o�/�/��u��$UI_PO�STYPE  ��%� 	�e�����QUICK?MEN  ��d������RESTOR�E 1ݏ%  ���,�>�b�m]����� ����Οq����(� :�ݟ^�p�������Q� ��ůׯI��$�6�H� Z���~�������ƿؿ {���� �2�D��Q� c�u�翰��������� ���.�@�R�d�߈� �߬߾���{υ���� s�%�N�`�r���9� �����������&�8� J�\�n��{������ ������"��FX j|��C���x���SCREր�?ۍu1�sc'�u2G3�G4G5G6G7�G8G��USER�).@T(IksTQ�4�5�6��7�8���NDO_CFG ޖ��  &� ��PD�ATE ���None V���SEUFRAM/E  ��&!�RTOL_ABRqT1/��H#ENBR/~C(GRP 1����Cz  A� �#�!��/�/�/�/�/B 6
??A*ՀUr(�A!a+MSK  hu%}1a+N.!%[��~2%��?��VIS�CAND_MAX�s5I�](�0FA?IL_IMGs0`����#}(�0IMR_EGNUMs7
�;�BSIZs3&����,CONTM�OUQ u4��|PE��c�� �@���"FR:\��? � M�C:\RC\LOGn�FB@� !�?��O�A�O_�z �MCV�O�C7UD1*VEX3[�Q`�qF�"ᖉ�`�(��=��͍_��Z�_�_�_�_�_�_ �_oo,o>oPoboto|�o�;PO64_9C9�B ��n6�eK CLIA�j�h�aV���lf@�g�o� �=	�hSZV�n�;���gWAI�o�4STAT �+B�@�O���z$����5J!2DWP  ��P G)�����a�;@'��2_J�MPERR 1�
  ��2345678901|� ������ď��ɏ�� ��B�5�f�Y�k���<�<N0MLOW{~�@��0�@_TIYH�'��0MPHASE'  %���3�SHIFTO21"x[
 <���?\� �;�a���q���Я�� ���ݯ��N�%�7� ��[�m�������ɿ� ٿ�8��!�n�E�����*	VSF[T1�cV�0M�ç �5�q� � �~�EA�  B8������ p������1���B ��ME$�u4�����a{~&%�J�M��x[�p�30��$xpTDINE#ND]H^8t�Or0U?��[J��S�ߏ���s5����Gy�	�߀,�������ߍ�RELE �s/q�XOjF~t�_ACTIV��x~8��
 A �;0}�<���RD�`���C!YBOX �X����v��p2���>�190.�0.��83��N��254�����`�� �q�?robot�ę�   pH<a�upc��� u��p��r����ZABC�#�-, u� �r�5X? Qcu������/�0//)/f/�Z;D�q���