��   9�A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����PASSNAME�_T   0 �$+ $~'WORD  ? �LEVEL  �$TI- OUT�T  &F/�d $SETU�PJPROGRA�MJINSTAL�LJY  $�CURR_O�UwSER�NUM��STPS_LOG�_P N��$�T��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD f� DV�IN!�$C� CRE��PARM:� T:DIAG:)�>LVCHK!FULLM0�Y{XT�CNTDސMENU!AU�TO, �$$�CL(   �S�����	��	�?VIRTUA� ���$DCS_CO�D@����� � W'_S  J*�! T&�Ar91&"!. 
 $���~-�/ �/�/�/�/�/�/?? 0?>?T?b?x?�?�?�?��?��`#SUP� `l+�?�?`#F�?�OFO��  �sLpA���O z ��� V�[t&�#�j�� mBO�O���G�O��XU 