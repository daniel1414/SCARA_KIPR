��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
GPCO�UPLED1 �$[PP_PRO?CES0 � ��1��UREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $,NO�/PS_SPI_oINDE��$D�X�SCREEN�_NAME ��SIGNj���&PK_FI�� 	$THK�Y�PANE7 � 	$DUMMWY12� �3��4�GRG_ST�R1 � $�TIT�$I��1&�$�$��$5&6&7&8
&9'0''�%P!'�%5'1?'1I'�1S'1]'2h"GS�BN_CFG1 � 8 $CN?V_JNT_* ��DATA_CMN�T�!$FLAG�SL*CHECK���AT_CEL�LSETUP � P� HOMEg_IO� %:3�MACROF2RE�PRO8�DRUN2CD�i2SMp5H �UTOBACKU�0 � �	DoEVIC#TIh��$DFD�S�T�0B 3$IN�TERVAL�D�ISP_UNITܻ�0_DO�6ER=R�9FR_Fa�{INGRES�!�Y0Q_�3t4C_CWA�4�12HGW~0z�$	Y $DB� �� COMqW�M�OJWH.
 \v�VE�1$F �A�$O��D�B~�CTMP1_F�E�2�G1_�3�B�2�GX_D�# �d $CARD�_EXIST��$FSSB_TY�PitAHKBD_YS�B�1AGN G�� $SLOT�_NUMZIQPR�EV��G �1_�EDIT1 �� h1G=H0S<?@f%$EPYO$OPc �0LETE_OKR{US�P_CRQ�$�4�VAZ0LACIwY1�R@Pk ��1w@MENP$D�V�Q�P��A���nQL*OUyR� ,lA�0V1AB�0~ OL]eR"2C�AM_;1 x��f$ATTR8�MP0ANN�@��IMG_HEIG�HQ�cWIDTH��VTC�U�0F�_ASPECQ;$M@EXP;�@�AX�f�CFT X $GR� ҷ S!1�@B`NF�LI�`t
UIR�Es3�tGITCH�~C�`N.0S�d_Ld�`�C�"�`EDkp*;tL0J*DS�0>0��zra�!hp;G0� � 
$WARNM'@f�+P� �s��pNST� CORyN��1FLTR�u�TRAT@0T�p  $ACC�1�
� ���ORI�	`!S<{RTq0_S��B�qHGI1� [ Tpu3I�8�TYVD+P*2 ��`v@� 1R*HED�cJ* ���2��U3��4��5��6��U7��8��9��qO�$ <� #p5x�s1v`O_M�@��C t 0E�v�NG��ABA � �c��YQ������@B������P�0X����x�p�P@yP�2� ����J�S_R��BC�J�L�2�JVP�CR���}@w��u�@MM�7CP_}0OF� 2 w @� RO_�̧��aIT8C��NOM_�0�1åq34 :�pPT �#�d��@xP��J}EX��G�0� .��p�
�$TF`��C$MDM3��TO�3&@U=0^�� �H�2J�C1{�E͡� vE`�uF�uF���ho@�a� 	P$@`�PU�3�f)�"��)�AX 1rDU�6�$AI�3BUFpV�o@�! |�plڶ�pPI��PZ�MY�Mf�̰i�}FZ�SIMQS� �/��A-������kw' Tp{zM��P��B�FACTqbGPEW6��Ҡ��v���MCc� �$�}1JB�p;�}1DE�CGڙ�G�i��a�� ě0CHNS_wEMP��$GO����+P_��q3�p�@Pۤ��TC��{r��q0 �s��a�/�� �B���!�	���JR!0��SE�GFR��Iv �aR��TjpN%S+�PV!F���ʹY��K��a1�)B���( 'j�Av�u�c t��aD�.0���*�LQ��D�SIZC������T��O�����aRSINF�����jq@��C��C����LW�8����x�CRCLuFCCCkpy�����N} ���bA�������d�*��DwIC��C���r���+ P��z�2EVT2�zFH_��Fp)Nt/�>�����H�1Q��!  ��@�Qx����U�kp �2 ��a��s�+���A|��S!x "� 4�4u2��tAR���`�CW�$LG�p��B@�1�Pr�P�t�aA?@�z�ϣ~0R�ӲM�E�`8�oC�RAs3�AZ����pb��OS�FC�b�`�`F�Mp�� �0��ADI S+�aV%��b�z��p E$�pRp�cV�S�P�L�a+QMP5�`Y8Cz��MeD�CU���aUS" $=�TIT�1�S�SG1���#�8��DBPXW�O! T#��$SqK��2�DBTm�TRLS$l�Q0T�Q��P`P�D�q�1L?AY_CAL�1�R^0o f7PL)A�Q��D'a�73a�7��	�)2!S%2?�PRj� 
*0���Sg& =�A$��S$ �*�L�9'�?�'�U�T(O�AS��PCS)#ODENE��*BO'Ӳ0�RE�pB+H ��Ou�&$L�C'$�3R��K2��LVO�_D~!U�ROSbrq�v�R����C�RIGGER�FP�A�S��6�ETUR�N�B�cMR_}�T�Ubp���@EWM$���GN=`���B�LA��TUܡ($=P�)$P s�*hP3a��C�TΣ@DO>���D�A���FGO_AWAY�B�MO"�a�!*0C�S_P,<aISt�� �� �s�S#�Q���Rw�cV���Qw2�VW��'dNT	V(��RV;����~���mgŃ��Jt��<@���SAFEڥ�f_�SV�bEXCLUtT��� ONL����cYfЀ�y�OTE�uHI_V} ��P�PLY_�q7�VRFY_b3���Rj L��_ -h@0��_�y�1� #tSG�  .�rŐ1P NQcQ� _q���;P���Vby|rsvANNU�N<@�$�tIDX�UR�c[P� �y�qi ��z�v��Ͱ�PI<B/���$F�r�$АO�TQP�A $DUMMY��&���&����*0t�U0 `  �HE�\����^r�cYRr SUFFI���Pa0��P�)�5#�6#�)1M�SW�U1 8��KgEYI��4�TM�A0��ځ3QՆINݱv��(2j P2 D��H7OST�0!��������������E�M&����*0SBLv� UL��3 Z���D�*0T�@S4� � $���USAMPa༥.�������V I�@��$SUB����;@c��8��3��SAV������������`�vP�$�@EC!	0YN_�B35 0��DIįt�PO\�M��#$�E�R_IB� �?ENC2_S�T!6X��2������  �cG���0 S72���1��A����8 � ��Ǜ��@PK��Dk!uq��AVERpҁ�����DSP�ܢPC?���26�\������VALU�HiE �M_�IP(îܣOPP� 5�T!H��ͫ��S` 4�.�FB�6d��~�� �5�SC?q���E�T�9ȂFULL_DU���qKP��0������OT�"�Q~PNOAUTOS:�$YĪ�Z� ����X�C��h�C�E26(1V�L� �;H *h�L � �����$P�� wc�ě1�Ʃ1��C���P���Ʋ���7��8�ɥ9��0����1��1���1	�1�1#�1�0�1=�1J�2X�2T����2��2	�2�U2#�20�2=�2Jڕ3X�3��3����3�	�3�3#�30�3*=�3J�4X�'���;SE�2< <8�Z����I��e�$�}��"qFE5P?PT= y,f��a? �PF�?i��e�i�E�Pq��aT�>F�$TP$!$VARI����7UP21p? 7���TD��s��p�������   ��BAC2@ T����$uP��*��Þ0� IFI@w�0�P� � )PB"�N�0P�TAt ;u�"�"pu STvt: �bt�@��l�6	sC2	 >0���S���/bF���FORCEUyPsr��FLUS�p�HfNn����bD_CM�PEv*�IN_t�e`�REM� F�a�a�0P�Te�KdN~��eEFF�j�PI�NJa�OVM�O{VA�TROV���DT	��DTMX,A��P*��0`M(xR#�0�CL*A_��u*�Pr�{_X�F�_T�+X��P%ASaD% ��(װ`�1`�&_APRQ�?LIMIT_�4�2� M��CL�tˑ�RIVW�*2EAmR�IOxPC�Pd���B�R�CMQP�*�b !GCLF�#�1DY�8} �q6�35T�%DG����0�5`�FS9St0��B P��1�A��`_�1�8�1�1��E�C�13 K5� F�GRA��gC���k�`W�ON<��"EBUGwctB�x#pC ��_E �D ��K� �/TERM�EE�EP�O�ORIS�@F�EcP�SM_�`���@�G�EA��TA�IHܙE���UP��Ig� -�Q��D|`|�C|PE$SEG#Zv�0EL�eUSE�PNFIzLRT�kAx,��DTF$UF�`O�$\��a�P/���Wi@T��t �cwNSTTPAT��<h��RPTHJKa-�E
�65MR<p&�WUw��&�Q�LQR<`�Y�qS�HFT��MQ�Q�X_�SHOR�*��F ��@$�GM`H�u O#VRq��q6`I`4�U� �aAYLO���"J�Iu2b��Q��oƸ�ERV���a�  6j�WnP�R~�E �eԌ�E Rb1Pp�AScYM|�p�MQWJ`W�� E���Qy�b0�U7tnPI��Uw�/�eaPo��`o�fgORnP�M�S�GRSMTfJg�GR��aC�q�PA|P��p=��K� � FT�OCFQ�P9`N $OP@/��#���N �!O�ڐRE
�RdS�QO����Re�R�UN�%�a�#e$PWR0IM@��bR_ ���=�.mR LVBH��_ADDR$�H_LENG�Rǁ����T�R� SO�M H�S���~�������	�SE!u����S:�MN�1N���p��F¹�O�L��8�3�3�=��ACROc�z�P$���[·a;�  �OUP���r_�I���q�q1�ѭʓ��ԙX!՘ Y1՘t!՘	�ԙл&E"IO���DϗA�xߕ9�gO $��<�p)_OFFb�;��PRM_Ò��H�TTP_[�HjP; (��OBJ�2���#$$�LE�S|���Q � �.��AB_�!T��椱S�p;x LV��K�R32@�HITCOmUBGE�LOہ磴!��@��"�Gf#�SS��HWD��SQjR�lpIN�CPU4BVISIO�����Ğ�
�������	� �IOLN�S� 0C�$SL�r@PU�T_�$@��P�V0� ʰ)F_AuS�2T $L  �� =a0U�@9`dQaٵ��䳊`HY#�0]�6É��UO�3U `"�{�$�5"M�5 Tƥ�R�P;@���`��T��µƊAUJe�V]���NEfgJO9G{W��DIS��1K��� �3W XХQqVv��P;�CTR�S�:�FLAGBB�LG�tX �� ���~aCLG_SIZ�����d �����FD��I�اؓ�׏ث@ �֎����	�d 	���	��	�@	�% SC�H_��R���aBg�NTє�Y��!E�2��p�J U}�}��p�L��|�DAU��E�A�����t���GHt�r���%�BOO�Zh A<�f0I�T2���@8�REC��SCRB�=�Dx:�����MARG� <18��0��a�%�	Sȣ$�W?�%���0��JGM��MNCH|z%�FNKEY���K��PRG��UF���g`��FWD��H]L	STP��V���mP������RS;	Hp��-�Cid6r0�.0s��	U|���r�Xb���P�E���G��`P�O�
.�M�F�OCU�RGEX.,�TUI��I��p�K|�V��V����A`B���p�A`�Nu��SANA%�FR��oVAILy�CLP1~uDCS_HIyD��
��O�X1�S�� ��S�V�IGAN��~�ӽ�\�T����_BUFF�1[j5�o`T�$��� ����B�P$��1\5�o`ܰ��c��pWOS1�%2�%3�!���_��0] � �ܩ�qEU�����IKDX�tP�bD�O� X��Q6ST|�R���YV�@1 \$EO6CO;�{�^6q68���1^ L��K� [@`�9`(��S���:������x��_ _ o�p�Ð��� C��@Cp�` �� C�LDP|�uTRQ�LI��Ft
�4I"DF�LGV�"@1VC�D)�VGr�LDVE@DVEORG
�qiB_�g��H
��d�D�ta A�M�@Dr1DVES�p�T4@I��@TVRCLMC%T�O�O7Y����MI��tb Ydy��!RQI�M��DSTB�0 ؓVO�XAXr |�X�\EXCES6���!vRM_��qc�0��Rt�V<��pd��V_A�Z��(k�_�X:@K�te \����n/�$MBs�LI��~�cREQUIR�b���l���hDEBUT��sQL�0M,�f�r�=��`����%RsQND���p�pgw�n�?�fsDC��IN�� ��p�,x' NV��ܖK�NA�cPS�T� h��LO�C�&RI���%EXvÀ�!�QsQOD�AQ,�i X��ON���MF\����v�9�2%��5�uk�0� w�FX�PIGG�� j �M��2!����3��4R �% ?3;�|�K�|�Z�G`E�ODATA{'��E��U��b"���NZ"k �t $MD��I���)Ɔ ф��фH��p�`Ѕ�X�҃AN�SWe�ф�!'хD�[�)�r��P��l -�PCU��V�X@�uRR2��m D��a���Rd$CA�LI�P"�G�w�2N��RIN��z�<u�'NTEڰ�"nI����°r��ڰ_N��o@Õޒi�oT۔bp�7DIVmVDH�Pݐ:��q� $V��+sv1$��$Z�"���� �"f�_�e�r�H �$BEL�T>��1ACCEL�!������IRC���P��t�T31h��$PS�P'BL�0 M�ʤ<C���������PATH������3ТZ��Q_�!U�2��8�R� C堌�_M=GP�$DDU���/�$FWh������q�����f�DE��P�PABNاROTSPEEH��!��4@�J��!��P���0�$USE_���P���O�SY��g�Q �B�YNyPAO��OsFF��MOUR�3NG�O�OL�L�INC.��q��u��Rxn�PP�RENCS������Rȡ���TŠIN�'2IТ���`R�V�ES�{���23_UyPI���LOWL!A� �4@���D� @�R{`���0��5bCΐ���MOS4 LdMO����PWPERCH   �OV��b� �!m�@1�^T@1�s�� hP�`�� V5�'`ѡ��L���Ig�����UP�Ӛ���TR�Kv�#2AYLOA A��$a1�Т@�5�p40��RTI(a|�40MO����R$b�@N��T��w�L���"f��DUM2,�S_BCKLSH_CТ ��B�A�u�'�Y�������6�x�aQCLAL�z ���Ar�`�CH�K4@+5SH�RTY@S��}%�A��_:3N6�_UM(`n�C{��c�SCL��ʰLM?T_J1_LS��P������E�����p������SPC��0;���	��PCsѦ�!H�0�`Y�q�C3P�2sXTc�g�CN_��N��i��SH ���V	�*3�Ň�=Т�2AC� y�SH:3�� g��ƝA���s�4�ѡ���c�PAx�l�_	Pw�[�_5@��8�V�04AH�ZK�JGG"M���OG[��TORQU��ON.�Q靰`wbLҠᝰ�_W��1�_A��G��M��UI�I�IM�F�p��JPQ2(�A_�VC"��0�T�RS"1Y.�P8m/�R`%JRKY,�"��&PDBL_SMth�RM)p_DLG�RGRV��$G��$M��!H_ �#�:�COS;`�8LN � ;;\%B4G�=9M�=9 !y:g<-!�%Z60L�ƾ!MYD1�8$2TH|*=�9THET0�NK23M�BA�E0[CBFCBA�C�Q��R,B$:AG�:AFSqBG�XBEGTSaʱC��qW4&�Dxg3�Gv3$DUH� Ih�Aw�x��R�F���Q9Q���v$NEd�AIF0Y�`R�E��$%��1A�5#U,W
581�LPH(eR��RS \%tSg5tSv5R�6�S(�Z�6%�VEXV:X7��]\VlZVy[V�[V��[V�[V�[V�YH�EX^Vdb\]�{hy[H��[H�[H�[H�[H*�YO6\OEXO�i[^UOlZOy[O�[O�[UO�[O�[O�6FR�'A�yg5�t8WSPBALANCE_�1��sLEo@H_�5S�P��X6�rg6�rv6PFULC�x��w��v5Ț1n}�UTOy_C�nT1T2G���2N*�z���g���@k���@ע����T���O����INSE9Gz�%�REV��%����DIF��1ol҇�1p�@OBȁ��#��MI��5��$?LCHWAR�����AB*y�$ME�CH0A�0>�D�Y�AX>�P��]�W(�<��q 
^������ROBV�CR�Ҡ�R=[��MSK_�pj�_s P R�_��AR��H�Ҕ��1����ԲҐ����Ґ&�I�N���MTCO�M_CD n�t � P�ڀ��$N'ORE��9���(�ou 8�GR��I�SD�@ABJ�$XYZ_DA9Q<���DEBU��M���U�v �p$�C;OD�� ��o��J�j�$BUF/INDX԰�����MORœw $1�U��-��v�F����ѣ�Gܢx �� $SIMUL�X�����$���OB�JE�p$�ADJUySB�5�AY_Io«�Dc����G�_F-IJ�=�T��� ������������Հt�P��D�FRI��׵T��RO���E�����OPWOܱ ɐy0��SY�SBU�PΠ$SO!P���#�'�U&�Հ�PRUN�M�PA��DL�H�!���_O�U�!A���r�$^��IMAG��ϐ��@P��IM����I�N� u£�RGOVCRḎ>°Ѐ�P����԰�@L_:����Lm� RB� �@�M��EDՠJ� 
��NpM.�������SL�pɐz x �$OVSL��S;DI��DEXqk� i�=!{��Ѕ�V���N�Ѵ{��Њӟך�ڷ�M�!E�_SsET�ɐ{ @����g���RI&���
B��_4A��	������ׁ@��  | HxϑI�J�ATUS��$TRC�@ǰˢND�BTMM�7�Ij����4��#�,�ɐ} DϐE~�k�A�`�EۂBᏱ
��B�EXEH�Z�ќ��{�b��~��АG�UP���$����XNN�m�=!p�L!p� �P�G&��!UB�6�g��6�
�JMP�WAI� P��N�L�O��1�F��#�$�RCVFAIL_C�1�Q�R��Q�Z��M� 𣕠���0R_{PL
�DBTBm��1�BWD��A�UM���IGe���m��� TNL� ����R���.�Ep�һ��!�DEFSPy� �� Lϐd�7 _8: H�HUNI��r��F ��R��^�� _L���P@���P�ȑ� ���F����Ѐ��p�N�pKET�}�r� P��ȑ� hW�?ARSIZE��l�h����S@�OR
�?FORMAT3���cCOJ����EMV�lUX�����PLI��ȑ� � $#�P_SW1I�-��AX����?AL_ ��E �A��B�,@C��Dnj�$E���u�C_��	� � �� ���qJ3x�@����TIA4�u5�6��MOM��@�����#�Be��AD�&�&�PU;@NR�J%�J%��DŔ�� A$PI�F�ޑ��$ �%�#�%�#�%=D�&�+ QD�DpсF���U�|��g�SPEED�`Gd*4f�7167f� ��16g3@8��O9��f�SAM�p맣417�3f�MOV���D�1@ƀ�E�4�E�17 1��42�������5n2��Hm��3IN2Ln �39HUK0Df�;J{HRD<{K�KGAMM�v�A>�$GET��Ƞ�L�D� �
b�LI�BR��I��$H�I��_��P��bVEĂXA^:P+VLW ]XVO\:Y|V+V�V������ $�PDCK�U�L�_�0�� �.B�m!E��W��T&�Yr ��$I�RS�D`��&����(�LE�`ޑ�Oh�)`�	E��ɐ�P��UR_SCR��a^���S_SAVE_DX�īe��NO�C� ���`�D��&�i� �)�iapz{p���& Ex@�q��0�B���5 G�2�+8!�;6��g8@�w�ucs�1��L.`Ŕ� ����!G�����c�w���`ζ�qW�`��$��0�N �d�R�qM��H�CLG��GM�aǒ� � �$PYr�$Ww�+�NGt��w� �u��u��u����@����@[L�nX� 	O�mZ��GQ�ŔG� pW�#�c�&��o�o#5��_)�� |Wи�`� �������`�ޗɖr�EQ��E OE����b�Ϡ���Pn��PM��QU�0� � 8� QCsOUa1�QTH���HOL��QHYSfES�1[�UEG�t�b� OM�  �1P4�U�UNI�J�� �O��)�� P�������a��GROG�j��2���O𤥥c�󠉠IN;FO(�� ��ث��
��1OI��{ (`SLEQ"6@D�5D�ܦ����DS������VPO�P�0#35QEMPNU�����AUT�a��COPAY�1�಼��`M���N������CT�� ��RGADJ(��2�X#�_$� '��'�W%�P%�]`'��:3�;�EX��YC���1@OՐ(����_NA�1!�S���i����M�� � ��p�PO�R��Ì&��SRV���)����DIT_p��� ��
��
�Tw�
�5�6�7�I8��1S�b�����OMC_Fe��p!L�a�a�;�Rq� ��/��җ#�0��k��7� ,`FL���ᦶ`YN{���Mp�C��PWR�����=���DELA �6mY�ADR�_j�QSKIP{%� i�����OŀNT�1�0*�P_����I� �`߂̐`��#`�3`� �n�kn�;�m�H�m��U�m�b�m�98a�Js2R.0��� 4� EX�@TQ��� �q���������jwRDCx�� ���
X��RF�E@AY��_�X�DRGEAR�_�@IO�t=bFLaG���EPC�εUM_���J2�TH2N�# � S1�UA�G�@T�P' �"���M��-�qI���4s!REF�1�1(�� l!�E�NAB� ��TPE 2`{� 8Wܠ�M �q�CL��R�w��
2'�-?Qc(u��3'��������4'��'9K]o��5'�������
�6'�!/3/E/W/(i/{/�7'��/�/��/�/�/�/�8'��?-???Q?c?u?�SWMSK(������ E�aMOTE���
��`/B`�L�q-CIO�UQEI�0��pPOW\`��� /���-������򿠨�ՈB$DSB_SIGN'a�q�����C��pS2�323E���$�DE?VICEUSKC�r>�rPARIT!�A_OPBIT�q��OWCONTR����q�0�rCUPM~�sUXTASK�S�Nq��P�DTATU��pS3`����u�e�_�pC��$�FREEFROMqS������GETA`.��UPD��AEbfS�PTP���� !>�8$USA����x�9h�{�ERIO��L�`ՐRY�U�B_�`��P�QQfWRK��?�<Dh�3fh��6F�RIEND�qg��$UF�U�p`TO�OLwfMYd�$�LENGTH_VTߤFIR��cM��SE�@�iUFINttrаARGIa�F�AITIi�gX�F�i�fG2�WG1`�� �Sr$wPR��sau�O_�@�P��xQ�RE���SU�ءT�C�N�=qyv �G(��]R���u��Q�A ��hzhZUz�ZU�t����{P�T�X T�P��L��TcH���hh�U�T�SG��W$X�)��r>�D����.��C�z�N�b��=$�v 2�!�-a�' 3i1?h.`21k2
��31k3?j���@i�����6{��s{��r$)V��bV�eV���vYr���O�[V{�@���hv3Ru�^pib��P5S��E�$���c��5$A8й�P!R)��u,�S���@����T�¯ 0�p�v���P�N�����!��P>p ��
�US^zA� �\�R���GA_�Š��Ny@A)XQ��Ag`L�ag�^p�THIC'a��8-����QTFE���>m�IF_CH'cp�aI_����6D�G1՘�٤*��h��`��_�JF�PRW�I���RVATF�� ��\�'�f`��)�DO��e)�COUW�C�A�XI�D�OFFS=EZ�TRIG�sz��,�)�#g���z�Hx����g�IGMA�P��a\���ȸORG�_UNEV#@Ͳ ��SD���d ӎ$����GR3OU[A�TOa�Q��DSP#�JOG�V�S8�_PV�3RO����U�mpEVKEPF��IR?�_�=pM �&��AP���E�������SYSv��B��;PG��BRKYr����b�\���������k�ADVQ�y�BS�OC�C@N�DU�MMY14��`S}V�DE_OP1S�SFSPD_OVR���C~�N�QÓOR\׶0N�P]�Fء�]�<�OV?�SF��a����F���Ac��As�؁a�BLCHD}L�RECOVM��P<�W�`M<��?�#RO1S�K�_a�_�� @���`VER�t�$OFS�`CV�@_bWDv� �rѰ��R��9�TR%Q|A�E_FDO�ƟMB_CM[A��B/�BLl�_¦�l�甁V�qDb�P����G���AM�Ú�yP��'��_M��>R��HC4�8$CA2���Ȱ>��8$HBK�Q��N�IO1e]�iAA�PPAQ�}�b���u���iB4�DVC_DB�c�񓡦B����A"��1��'���3��-�/ATIO�@��FP�M�UDc1�HFCAB H�0bFs�p�p��Ea�<�_BP��SUBCPUk�I�S%��@�� ��P�s�,���B��?$HW_C!���i��x�A'q\�l$�UNIT��l�A�T}����I�CYC=L��NECA#���FLTR_2_F�IҤ�H)�FEaLPxU˲���_SCTosF_�F��
v�
�FS�A���CHA�Ja^���3R�RS�D1�B ё�l�i@_T��PRO ~�)PKEM�0_���8��3� �<�*%D�I�P��RAILAiC��rM��LO��c+�i���-��-V'�PR��S{q�0ҕ!C���@	&�FUsNC�³�RIN�p`Z�+`? �$(QRA� mr 9��#��G��#gWAR�:�BLuq��'4A;88D�A���!I835LD@�PA�A�q3h��!��q3TI���5�β�pgRIA�Q�BAF� P�A���1��5��T����EMJ�I1Q��D�F_�`�ӨQ��LM�t�FA�`HRDY4d�P�`RSoq+`|Q0EMULSE�`x���E� ���I�����$]a-$�Q$�Q�,���� x��EaG���AРAAR�2)�09mb�E50��wAXE&�ROB#��W�ac�_�M�SY����Ae�VSWWR�ذ�M12�� STR�"Ņ�d�h�E� !	CUq#��lqBhP3�oV��)��OT�Pv� 	$�ARYg�ЦR_!�`	T�FI���j�$LINK(�1w��Q�_eS3��CU��RXYZ@Q��[��	co��Q�RJ�X�PB!��"Kd0�
 � LcFIeg`3�D�9Ԫ$<�_JN�p"�e��SA�OP_~T2�[53�NqTB�aNB2�bC9��DUQ�BV=6r%TURNb����u�Q�!h�?�gFL�)���B�@+pekZ7�3�I� 1�nPKH�M��BV8r%����c�ORQ&�!�# mX�C�����갦��up��.�<��tOVE�q��Mj�tC�zC��B�W�Fq�� � ��� j�0���qw�P� ���	��q���zC��L5��!ERM��!	v"!E8P���#؄A���id�%"�WP1MP1AX�bP1��&!�Q2� 2!>�\A>���=��`=� p=�ep=��p=��@=� JQ=�@:�@J�@Z� @j�@z�@��@���@��@��ב˙DEBU�$�!�1($�{�P��R�g� � AB�P'N�[��sVְ� 
����Ϥ��Ϥ aڧ$aڧ�aڧqڧ eqڧ�qڧ�A�4�`�2\�RLcLABbb�u� ���1s  ��ER�9P �� $8`� A�!��POB�FЉ�P��ލ�_MRA��� �d O0T<�\�EcRR:�2�0TY��aIA�Vb`,���TOQ+�i�L�@,�7R����� C�A � p�T�P��< _V1ْ.�V�2#cą2\�2k�ȱ��op�8ˠȱu�$W��j6�V�A���$�@"�0,���6�Q�	�@�HELL_CFG��A� 5e Bo_BAS��SR��\p�� �CS�T�1�1��%�22�U32�42�52�62�e72�82��RO ��8��P,`NLzA�cAqB��H �ACK�� >�i���`�`G@���7_PUr�CO�@��OU��P0�W!���3�7LTPX�_KcAR���RE���&@P W1�0QUE�� �p9CCST?OPI_AL������PU#�Д���PSE�M���M���T�Y��SO��W�DI�����}�L�1_T}M�MANRQ���PEZV�$KEYSWITCHU#�8��CHE9BE�AT!�!E�@LE(�$f�U4�F��5�|K��O_HOM�0�O�#REF�pPR��!)�AUP��C��Op�0ECOư_1`_IOCM�d����Q����g�@� �D�Q� U۲{�M�w2Q��p�cFORC��3 �p��OM>�@ � @���3*�U[SP�@1��$��@3�4�1��N�PX_AS�¼ �0�ADD' h��$SIZ�$VsAR2�D@TIP��)�� Ah�аJ� � �� �BS��AyC��%FRIFa���Se�w	��NFp�@Џ@� x�SI�TEFsj"es�SGL}T�R7p&�A���#P~STM�TJ�P�@;VBW<�pSHOW�R���SV
@�D��; �ԱA005pЁ  "� '� '� '� �'5)6)7)8
)9)A)�@'v  'V�	&r`'F(JP �()�P�(,)#`�(F)@p�(`)�p�(z)1�)U1�)1�)1�)1�)U1�)2)2)2)U2,)29)2F)2S)U2`)2m)2z)2�)U2�)2�)2�)2�)U2�)3)3)3)U3,)39)3F)3S)U3`)3m)3z)3�)U3�)3�)3�)3�)U3�)4uI4)4)U4,)49)4F)4S)U4`)4m)4z)4�)U4�)4�)4�)4�)U4�)5uI5)5)U5,)59)5F)5S)U5`)5m)5z)5�)U5�)5�)5�)5�)U5�)6uI6)6)U6,)69)6F)6S)U6`)6m)6z)6�)U6�)6�)6�)6�)U6�)7uI7)7)U7,)79)7F)7S)U7`)7m)7z)7�)U7�)7�)7�)7�)]7�$Q�Pd��UPD��  ����)и�YSL}O��� � �`��Q��TA��8�����ALU���Ц�CUT��F��IgD_L��HI��IV$FILE_��?�+�$����S�A��� hҰk�E_BLCKh�x��>��D_CPU���  ��� �B�T���q�	��R �G�
PWll�� �LA1�S������RUN u������8�u�?����?�� �T?�A�CC��X ;-$f�LEN��s����f�����I�J�L�OW_AXIh�F)1f�,�2��M��	�G�_��I��Y�8�թGTORn�f��D��<ܣ\LACE��Y�pf�ٳY��_MA� p��3�	�3�TCV:�[�	�T�\�{�q�| ������	���J���ŉMĴ�J9�����	�r�2�Ц��������ΠJK�VKо�#���#�3�J0l8�'�JJ/�JJ7�AAL'�]�/�]�W�e4X�5��{�N1��P��M�I�ڤLӠ_����b���� `u�GROU����}Bd NFLIC���REQUIRE��EBU��b�Ŷ��2�c�	�a�� ��� \APKPR�C �ܠ
a�;EN\�CLO��lهS_M`������
�a��� �F M�C6�{�����_MGV��C�l��؎�5����BRK��NOL������R�_LI��������J��P _��/��7��{��D���6L�O�8���b�?��� �ҍ�z��燡��PATH�������ᒨh��� $��ͰCN���CA �]���INFe�UC٠��%�C��UM.�Y��4���Ez�P���P�7�P�AYLOA�J2=L��R_ANE���L���������R_F2LSHRC��LO��$���2���>2�ACRL_�"�� �����H�b��$H��CFLEX�_�`�Je�� :r���	�t���`��	�������F1� ��ïկ�����E'�9�K�]�o��� �������$��гĀ#(ؿ�����TR'�X ˲�`H ��%�&�8�J�\�`� i�W�{ńϖϨϺə�}J��� � ��0����ʁ��AT�6ðELt �5صJ����JE��C�TR�TN"F��6	�HAND_V�B�_����� $f F2�֋���SWF������O $$M���R�Ӏ�H�ѕL��E:�FA@�������I��A��݀��A��A	��@��T����D��D	�P��G	�qYST��yQ��yQN�DY �Z��� �D�E��)��������@���H$� � �PT� ]�f�o�x����}3>�� {@`��n�xvf��o�ASYM������Ͱ����_SH��#�=�'��dLHG�Y�k�}���J���G��gs]y��_�VI/C�x�ӵpV_UNI���t�#��J��re�r���t�� �t�ð	G�(:$j��#PXW��AЙH��N��EB��E�N/@��DI	�W#OƷ� ��Й����) � �BI�aA;��� �吂��U��0`�瑾n�� � ]AM�E\?0�g���T��PTpi0��5������K�,p:�U�I�T�Kp�� $DU�MMY1�!$P�S_RF�   �����͑LA��Y�PV#��=�$GLB_T~@��ŕ5���p`�CAӁ� XIЬ	נ�STȱ�S�BR��M21_V�ɲ8$SV_ERb��O��#�CLߐ��AuO炔��0O�� � D fĐOB���3LO��f�S�y�ÐS�p�1S;YSS�ADR�1���5�TCH�@ �� ,f L���W_N�A
����y5S�R>��l  }J�J���F��B�� �G���I���ID���D� ��D���V�p�KYV��� bu���ݻ�������);Mt��XSCR�Ei�W��E@�ST��F�}��a�Ǥ���0_�0AV�� TI�&����1%��ࠬ���1�����O�PIS�1�����;UEЄ� ���SG��1RSM_�����UNEXCE1P��ј�S_ߑ���7��&�9�T���C�OU\ғ� 1-֤�UE��؂6��y�PROGM@F�L�1$CU&�P�O�>��I_�H>�� � 8E��_HE_������?RY ?�0���p������OUS� � @��D�_$BUTT/�R��>��COLUM0���s�SERV�3��P�ANE�0V���NTpGEUA|�F��~ʡ)$HELP��^�bETER5�)�� E���Oq��30��;0���M`��U`��]`��IN��-�TpNp��0��131� ��i�LN��� ��0���_����$H_�0TEX�3j�^񼪑~$RELV"DP��~Ӑ�b���Ms�?,��p��4�򪑥#���USRVIE�WV�� <���U:"�]@NFI�0���FOCUA���PR�I�`m��h� T�RIP��m�U9N��Є� �`/���WARN����S�RTOL��&�tRs�O�cORNs'RAUW�vT�	����VI�υ�� $��PATH����CACHV#LsOG��LIM�r��S��BR'HOS�TǢ!���R�|�OBOTƣ#IM� ��S���0r��������VCPU_AVAIL��V�EX�!�aN���} ~�Ma�Ua�]a� ����ƀ$B?ACKLAS� �!��$"W��  ��C�T%s�@$TOO�LǤ$�_JMPΤ� ���$�SS�v4��VSHsIF`у�PB����ǤЇ�Rk(�O�SUR�3W�RA#DI�$��_���%��м1�ぺ��$LU��q$OUTPU�T_BM��IM����b� }p���#TI�L�'SCO�"�#C ���$N�&N�'N6@N7N#8���u%(=,�2�TQ"�`rЄ�<��DJUr|U��P�WAIT����<��:%0NE�~��YBOW� ?�� $����v��SB"ITPEo�NEC/,B@D(D�PJǐp�Rv hE(�#H=@�0�B�E/�M�K T���"y�� An�!ӻOP�
MAS��_�DOآ�qT��D�]����C��RDEgLAY��SJO� "X֡�c'T�3��`� 0��,l�y�Y_R�y�wR�#ƢA�?� ��ZABC�� ��R���
  �$$C|�X����Q𘐎��P�PVIRT8�_�PABS�!���1 �U�� <  �Q(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П������*�<�K�`�AGXLM�0���Q�c7  �]�INf�x��\�PRE�Nk������LARMRE?COV �Y������@F �U/�QdK�� "�4�F�T���w�����<����, 
#o忶W�NGu k	? A   �,˾`PPLICu�?��U����Handling�Tool m� �
V7.70P/�36+��
��_3SWr�F0���� 43�ˊ�yϋ7DA7�철�
f��rm�N�one����O�հ�P�T���.�RAP_+�V��R�:v�7�UTO�RX �l���n�HGAPO�N�Pe� an�U' Dw 1�� ���������T�n�� Q �1�  �0��
����	7�H嵡]���R�R �a�,�H��B�HTTHKYV� �R�+�=�O������ 3����!�?�E�W�i� {�����������/�� ;ASew� ����+� 7=Oas��� ��'/�//3/9/ K/]/o/�/�/�/�/�/ #?�/�/?/?5?G?Y? k?}?�?�?�?�?O�? �?O+O1OCOUOgOyO �O�O�O�O_�O�O	_ '_-_?_Q_c_u_�_�_ �_�_o�_�_o#o)o ;oMo_oqo�o�o�o�o �o�o%7I [m���������!�[���TO��C�U�DO_CL�EAN��5Ի�NM  	�Կ���+�=�O���_DSP�DRYR��HIa��@����ϟ�� ��)�;�M�_�q�������MAX@���[����׳�X�����҂�>7�PLUGG�У�\��S�PRCt�B�E�������O��}�5�SEGF{�K Y�k�v������Ͽ�p��=�p�LAP�� ��o�Y�k�}Ϗϡϳ� ����������1�v�TOTALզ��v�_USENU����� ���ߎ���RG_�STRING 1�s�
�M�l�S3�
��_I�TEM1��  n 3������"�4�F�X� j�|���������������0�B�I�/O SIGNA�L��Tryout Mode���Inp��Sim�ulated���Out��OV�ERR�� = 1�00��In c�ycl����Prog Abor�����~�Statu�s��	Heart�beat��MH� FaulAler%	U�CUg�y������ ���۞����6 HZl~���� ���/ /2/D/V/8h/z/�WORy��� �!&�/�/�/�/?"? 4?F?X?j?|?�?�?�?��?�?�?�?OO0NPO��V@�+?OyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_p�_�_�_QBDEVYN �PmO�_!o3oEoWoio {o�o�o�o�o�o�o�o�/ASewPALT�q�/x ����� �2�D� V�h�z�������ԏp���
��GRI�� ��B���j�|����� ��ğ֟�����0� B�T�f�x�������0�j�R�Z���� � 2�D�V�h�z������� ¿Կ���
��.�@�<R�ԯPREG�~�� ��dϲ���������� �0�B�T�f�xߊߜ������������X��$�ARG_� D ?�	���9���  	�$X�	[M�]�M��X�n�,�SBN�_CONFIG S9�������CII_SAVE  X����,��TCELLSET�UP 9�%  OME_IOX��X�%MOV_H8����REP�S��&�UTOBACK�����F�RA:\x� XZ�x���'`��x�\��l�INI�px����l�MESS�AG������A���ODE_D����#�O�P2l�PAUS�VA!�9� ((O<����� ���(^�L�p��ej@TSK  u�����o�UPDT) ��d� ?WSM_CF��8���%�+!�GRP 2
5+� L�B��A�#�XoSCRD/!15+' �������/ �/�/??(?�����/ p?�?�?�?�?�?5?�? Y?O$O6OHOZOlO�?�O(�r�GROUN� S�CUP_NA��8�	r��F_�ED��15+
 ��%-BCKEDT-�O0�%_I_�� ���-r�_x�eo�o�x���UA2r_/��_�_�R�o��iU�_&o�_�_ED3 o�_�o�_n_o�o9oKoED4�oro'�o�nn�o�oED5 ^�:n����ED6��o���nK���%�7�ED7 ��^����n�Z�ɏۏED8J�*_��N_�m����m��ED!9�[�ʟm7����#�CR_��� �7�ٯD���ū�@�@?NO_DEL�O�B�GE_UNUSE��O�DLAL_OU�T ��R�AW?D_ABOR����AݰITR_RT�N����NONS�i ����CAM�_PARAM 1�9�#
 8
�SONY XC-�56 23456�7890H �~��@���?��( АZ����yŀ��\�HR5po�������R57����Aff��\�L� ^�Z��ߔ�o߸��ߥ� �� ���$�6��Z�l��a�CE_RIA_UI(%;�F�!�{�x� ��_�LIS$�c%����@<��F@�GP �1Ż����OK�]�o�.�C* Y ����C1��9��@��G���CP CU]��d��l��s��QR������[��m���v���������W C���& ��G��;�HEנONF�I���@G_PR/I 1Ż��T ������� ��CHKPAUS�� 1I� , �BTfx��� ����//,/>/�P/b/t/�/O������8�!_MOR���� ��@2C�3�������" 	 ���/;�/.?? R?\5�"����-=�ֱ?99��3�@K(�4��<P������a�-8��?OO�J
�?KO�'ưS��"��:O��i`��P�DB� �-+�)
�mc:cpmid�bg�Od��C:� � �PP���Ep��O-_�CP�7@�
7@�V�@�Oq_<Z+�.��.��S[_,�_=Y�,�F,���bUYg�_o�\�װ�S[f�_KoAMo�J?DEF ch��)�B:`buf.txtqo�Mro�0����'�	�A��1=�L���jMC�#��-,���>ss�$��-�r���Cz  �BHF3Cs7 C����C�M�F���iDP�E�~�WJI0D��tE�qaEp�IJ$�3H�HƷ��{G��G��GG����N[5K~�w)L��XWI>���{,�O�fu7���4�),�,�.*װ�,�,��@�u��K�x6�q�* ��* e�D�n��pE�WLI0EX�E�Q�EJP F��E�F� G���}F^F E��� FB� H�,- Ge��H�3Y�WI?��p�?33 ��%WD1n6��"��5Y��\2���A�1WDq<#�
 �O+�)�Zj�b�RSMOFS��ؐn6��iT1� DEg  �?DR 
�v,�;�&�  @��:��nTEST�bo�8�R��!�/3�nvMC+�A�WJq� [�Q�rq�C�pB1 Jw�Cy�@T�6���T�FPROG C%ź��ů��I����𦶠喤KEY_�TBL  �6Q��!� �	
��� !"#$%&�'()*+,-.�/01g�:;<=�>?@ABC�`G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~��������������������������������������������������������������������������������͓���������������������������������耇������������������������LC�K�X	���STA�T*��_AUTO�_D����G_�INDT_ENBK�b�"R��i�[�T2�Ϟ\STOP���"T{RL��LETE�����_SCREE�N "�k�csc��U��MM�ENU 1""�  <����|� WE[߅ߺ�V��߽��� ����,���b�9�K� q���������� ����%�^�5�G���k� }������������� H1~Ug�� �����2	 AzQc���� ���.///d/;/ M/�/q/�/�/�/�/�/ ?�/?N?%?7?]?�? m??�?�?�?O�?�?�OJO!O3O�OWi;�_?MANUAL�Ϟ�oDBCO��RI�P|�4�DBNUM�`��<q*�
�APXWORK 1#"�ޟ+_=_L�^_p_�[��ATB_�� $�"��ipT�A_AW�AY�C
�GCP� *�=���V_AL�@M��R�BY���*���H_�` 1����/ , 
^7�6�PBoo�f�PM��Ij���\@��cONTImM��*���f�i
�$cMOTN�END�#dREC�ORD 1+"�8er9�Q�O�Oq= 6��R{���Hx� �O�s(�:�L�� �������ʏ܏�  ���$���H���l�~� �����Ɵ5��Y��  �2�D���h�ן���� ��¯ԯ�U�
�y�� ��R�d�v�������� ��?�����*ϙ�N� 9�Gτϧ`�^�ϼ��� =�������(ߗϩ�^� p��ϔ�����9�K�  ���!�H��l��� �ߢ��K�a���Y���}��D�V�h���RTOLERENC�TsB�b�PL���@�CS_CFG �,0k�gdMC�:\��L%04dO.CSVi��Pc����cA CH z�Poo�n"W^m�c���RC_OUT �-�[=`�o��S�GN .�Ur���#�05-�JUN-20 1�3:15 �Q�25-MAY�1�:00 af P�X��n ��pa�m��P�JP�{VE�RSION ��
V2.0.�11�kEFLOG�IC 1/�[ 	tH�P��P���PROG_ENqB�_r�ULS�g� �V�_WRS�TJN�`�Fr�TE�MO_OPT_S�L ?	�Uac
 	R575�cVO 74T)6U(7U'#50y(t"2U$tH��/z2$TO  �>-�/{V_�`E�X�Gdu3PA�TH A�
A�\�/]?o?�kICTZ	aF�P00g�T>dceg��1�STBF_TTS��h�I�3U�Cda�6��@MAU ��bMKSW��10i�<�l� ��2�Z!�mO|3 bO�O�O�O�O�O�O_�tSBL_FAU�L� 3�_�cQGP�MSK��bTDI�A��4�=�d`���a1234567890�Wc|6P�/�_�_�_�_o#o 5oGoYoko}o�o�o�o��o�o�o\SpPf_ *��OR*�?%�P Bhz����� ��
��.�@�R�d�8v�H|��UMP4!Y3 )^��TRNBKS���ĀPME�5ЏY�_TEMP��ÈÓ3��D3����UN�I.��YN_BR�K 5����EMGDI_STA%��W�NC2_SC/R 6G��_�� ��͟ߟ�f����0�0B���~�e�17��;�������¯,R|�d�8G��a����� ��N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶�0�� ����@$<��)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ����������� �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/��/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgO�/�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo �Oqo�o�o�o�o�o�o �o%7I[m ������� �!�[oE�W�i�{��� ����ÏՏ����� /�A�S�e�w����������קETMODE� 197�v�� '�� �W�R�ROR_PROG7 %�%���X��'�TABLE  �A�������њ�RRSEV_NU�M ��  ����)�_AU�TO_ENB  q#��j�_NO�� :�
���  *�F��F��F��F���+E�_�q����HIS�h����_ALM 1;.� ���F�F�+�� ��$�6�H��Zψ�_�%�  ��D����ېTC�P_VER !��!F�j�$EXTLOG_REQ��s����SIZ��~��TOL  h�{Dz���A ��_BWD�5��a��	�_DIO� <7��	�h��k�STEPw߉�ې��_OP_DO��4��(�FACTORY�_TUN��d��E�ATURE =�7�a��H�andlingT�ool 7� DE�R Engl�ish Dict�ionary=�7� (RAA �VisS� Mas�ter0�>�
T�Ea�nalog �I/O7�>�p1�
a�uto So�ftware U�pdate�� "�`��matic �Backup;�d�
!��gr�ound Edi�ts�  25L�Cameraz��F�� "Lo���ell��>�L, �P��ommj�sh��8�h600%�c9o����uct%����pane6� DI�FD�'�tyle �select�-� `�Con��j�o�nitor<�B�H���tr5�Reli�ab�� �(R-�Diagnos���:�y�Dual� Check S�afety UI�F��Enhanc�ed Rob S�erv��q (V��User sFr���T_iE��xt. DIO V��fi�� Z�\=wend Err��=L��  pr�[�r��C  P���EN�FCTN M�enu��v����.�fd� TP In�p�fac�  
�v�G��pl�k E�xc	 g5t��High-Spe �Ski��  Pa�r\�H��G mmuwnic��ons��7\apur� p�~��t\h8��^�conn��2�{ !D�Incr� �strZ�i�<�M-�6< KAREL �Cmd. L� u�a���8sRunw-Ti4 Env=�(mqz m�+��s���S/W=�"y��License���' a���ogBook(Syo��m):��"M�ACROs,�/_Offse��f��b�HG R��M1?��MechStop� Prot��d �5
$�MieS�hif��9�B6SD�Mix ���7��y�Mode Swoitch��Mo��*��.& �M�&���g' 65�ulti-T� ����Z��Pos��Regi�o�  ! 7P>r�t Funb>��6iB/1��Nu!m ��dx�P`�31>2  Adju:��/2HSM7Z* o<Y�i8tatu1<�wAD RDM�otN�scoveW� #��3��uest 867�.�9oG � �SNPX b����Z#�LibrV�;�rt IE,� S$@��.�0�� �s i?n VCCM9��0�� ��!9�3���/I� 710~< TMILIB�MpJ0,@� �Acc�����C/2@�TPTyX"+QTeln ��Lq3�%|(PC�Unexcep�t motn�� �0�0,	7�\m72f�+4�f�K�  h64aVSP CSXC9�@(Px�U["3� RIN�sWe'50,D���Rvr�	menXS@� �QiP^ a0x��3fGrid�1�play F O``�fp@��vVM-�@A(B201 f`�2� ORD|�s�cii��load�3�41%�lJ�i�GGuar�dP�mP���k7�b]aPatv�& 0N"Cyc��0ori���`i�C00Data�@qug�c�3[,`�37FRLOAam�5<�~�3HMI De�2�(�1oc644�0P�C�sePassw!o�aA)qp�1p���\{-+PvenjCT����YELLOW� BO�I t�"A;rcV0vis���%����Weld� c�ial�$   5 �et�OpA ;�g41\\�5a 2��a��po)@`@�a�T1���50.2HT̰ @ xy�R:�82���`g�P��xp��� 12�AJPN �ARCPSU P�R\A�TEh0OL�wpSupg�fil�5p�Q��^ l�cro�6 "T�`�3E�Ldx�!��SSwpe�etex^$ J3ֳQSo�t� ss�ag�% T�eBP�� ] !9M�Virt���39�V h	`stgdpn6��ro� �SHAD�pMOV�E TF MOS �O � Dge�t_var fa�ils ��ߐ  Ȫ D��E��� Hold Bustd�CVIS UPD�ATE IR��C?HMA 62�q��WELDT�@S �) "���: R�741-�ou
�b���m BACK�GROUND E�DIT Ò m4�1�0REPTCD� CAN CRASH FRVRT�O�Cra.�s 2�-D��r �0r�$FNO NO�T RE��RED� � PCVl�J�O�P QUICK��OP FLEN/ .pc�c����TIMQV3 ld�m�PFPLN: �燹 pl 2���F�MD DEVIC�E ASSERT WIT iC���sANġACCE_SS M �aŀo1Qui��<!좝C"�USBU@- t� & remov���<�2� SMB �NULApܡ��FI�XW��HIN͑O�L2�MO OPT>t�PPOSTwp���D��- � �Ad�d��ad. 	�io֬�$P:�Wu`.$ZѠO��IN��M���CP:fix C�PMO-046 _issue�tJСsO-|�2�130����SET VAR?IABLESΐ�$�O�3D m�"vi�ew da`PWe�a�80b. of �FD ��u)��x� OS-1�p� hG s v�D�5t��;s ��lo �(�� WAx��"3 C�NT0 T�S$I�m�Z#ca��PS?POT:Wh�p��ns�STY܄At��pt�do GE�T_l���VMGRw LO�0REA�p	C��M`P�@ Y�|��0�ELECT���L��ING IM'PR N���Rɰ̐�sPROGRAM��RIPE:ST�ARTU�@AIN�-��D��QASCIyI�d�OF L����!`PPTTB: mN��MLKdme�4ڃ�:�moW�al�l��R� Nu�Qr�� Ang���`d���tho�n[� ch >`ܐ�r R2wtoun�H85@�iRCalA�"S'ign�0�pI,A��Thresh12�3�#.c�Hڰ : MSG_P�ю�per �ࠡ��A�zero5P� A�g  J�!O�Imr �� 2D�0rc i{mm�`SOME��s�ON������0S�REG:�^5� �LB A9�KAN�JIH�no��`c�	��n dq�� �-1o��INIS�ITALIZAT1I��we��0= dr\  f��aP����minim90r�ec 1lc0�:�?!blem��ro���L�<3a i� 0�9 ��b�d�w-� 8ݡ�0�w uHQm@[se�4SY�M��0s���QЧ 090�Wklu� E;BRe���jձ4�1���m ����Par�r@ G�B�ox fo TMyE�ːRWRI<����SY��\k��F�/�up��de-rela2Qd��#5��betwe�pIN�D��GigE s�nap�us5�s�po V�TPD���DOs�ġHAN�DL �`�Q�i�Dz��n�0 f.v����Boperab;il�` tmCQ��': H5@�`l��L�
! ��m@p�h�s UIFL�P�O>�FA����ΑV�7.��CGT��p�i�AsM�5pj�)@U���ine-Rem�arkO@0 RM�-�$ÔPATH {SA̐LOOS��ܓv�`fig�GLGA  �0%���p���J� ki q�the�r�A� Tr�`iEn�DW����2�7��� X�е���8`n&;� C� ��:  6��d� y* it 3w5\k�Pay�a�[2]_�D1: ug�s> dowD2�	SDISp�1�EM�CHK EXCEy ֠�$MF +  ��h�"�P��Վ�B0 ce1Ȣ��#me�� �c� !�?��bP�� BUG���yB
�@DŠP�ET��V0�0�T93~X�XPANSI)��DIG��O  �H5�P�CCRG� ENCCEMEkNT`�Mm�K 1�A�H GUNCHG OA�1Tڐ���
�Sg\d���10ORYLEAK�������LC WR�DN R��O�`j95`PO�SPEްC}G�V ont���VM����W��@`GRI,@A�7��� �PMC ETH�0�i�SUذ>� H5y7�P0PENS!��N���ː RE �(i�ROW<�³R�MV ADD  1II�=p��DC^ q��T3 ALAӀ ���m��VGN E�ARLY>���f n�� ��衸E�ALAYH7u�СPDg�ˀH1S=S8�OUCH��D���Fh�����PCDEoRROR*PDE��� WRO��CUR�S�PٰIp@N gxҰ�?Q-158Kw9a���SR �ġ9U3��\aptp��
@T�RF@�R�\`��UB�U �`��#RB��0SY RUNN̤��`10�ఱBR7KCT@qROq�Ԁ���CDAX��Djj�EISSUcހ\�\�D��TSI�aK�t�XM�IPSAFE�TY CDECK "M6���dѤр[`S U�)��4}P@QT�WD��E�'QINV��D ZO����a�xsb_aBDUAL@(|�'QòF��E�4l��6��P`NDEX� F�P�U���SUFrPk�Lbѳ�RRV�O117 Ay�Tp��챤 ��FAL�B�TP247���P�?q�EHIG�PCC� n��0�ESNPXV*PMM�Q ��)!SQ�"V��8T�bDC�B�DETEC��ds!Sˀ�BRU/b63�<��s� 02"�t�s$�'�!h� Z�T�7pSA��"e���߆��,@����߉ـ�0�
աx��ق�cscr��ـ �dctrldA.؁���fّ��!���fـ*��W878��-�% ��/� rm��
�Q�mR��78�RIـA�̑ (��~��Q .����ao�ـ\��a@:P���a��I��ta O3 "K:����<��#�o��tp؁ "PLCF"E!�ـ�plcf���ـ-���mai�ـN�F��ovc���ـt��/�ـ������􁢐r�674��Shape GenwـEI��R,���ـT�ь�V� (5�ـ��II���� �+��ـl�֟�sga 4P� �4j�I�r6ـŲ5�=�5ѺI���ets�6� " PC���n=ga�GCREѿ|�85��@�DATj����5ŝ�t.!��5�a�񯜳A�gtpadxb���Y�tput��@����ñ��2ـ`��5Ĺ�����sl�v�q� 7�hexy���4�����2�keyy�ـ"�pm������3us9ߜ�gcـ�����+�H�a�j�921��pl.Colly󔱾�r�В1N��ڕr� ({�ـip���r��'����8�7=�7���tp~�� "TCLSj�<|���clsk��D�:��s�kck��� )�U������r�H����71a�- KAR�EL Use S=p�PFCTNj��a7��a�a��� (�� ѡ�� �ـ��ٹ�6��8=�8"   ��ـ 0S�(�V�   lm� 6�99�~ F�|)vmcclmf�CLMl��`��60v3et���LM:��檡sp]��mc_mot���ـy���suX��p60���joiT�xJ��_logH��trc��ve%�� �����~g�finder���Center F8b!��M�520����lg��  (m)r,���fi��1��a#�z�� �ـJ��$t�q� "FNDR�����$etguid@�UID�ـ
?�1��E7�q1nufl�6 �ـ>_z#ѯ7A�x��(�2#���$fndrp����c$��tcpS$�]�CP M� H�3�ـ517��g�38 �vC�gD�*Y=�F�| Ց� ^ ���Ct	mgA4�P��O�CG1�ՑO7�Y��8�Et!m �?�Wـe�?�C�Rex�ے���Z8��ڔXprm؁�_|�D�_vars�_ Z$M���Vh@����`��gG��ma�w�Gr�oup�@sk E?xchang{@ـ�ÖMASK H5~�H593 Ha��H5���`6�`58J�a9�a8�B�a4q�2���b(�o#
k��/�غ`hp8�0Y0`/_цt�qTASKY_��r��pz�h�Z�m�@��������SDis�playIm��v�{Gـʑ8�OJq(�P%���@a���a��� ـlqvl? "DQVL�t���q�����Ϧ�y��|���1avrdq֏4ᩅsim���0��#st��o��d���������v�0Z樁����"v�Easy N�ormal Ut�il(in4�|+1?1 J553��a�Dc���(���0��)�M��<�O�<� k986�TA8��#�4�� "NOR�
��1�_���|�su��.������7����a!g�y! me'nuu��g#M���މ�R577� 90� ̒J989��4�9�L�A0�(�ity�E�A�,�P�m&&��mh8��"8 2��܄����C8_Sշ��n "MHMN �r%.Ը%���ͯ�s� ���i�Ը-at�Х_��������ֶ��tm��?мz�1����Q�2ȭϿ�z�3zos�od3st��
�mn�O^��ensu�Lm���hRaL�߃��huserp�a����c~���Ը5�ɯ��<���oper���X>Ըdetbo`Ý~  ��LUA���������dspweb ���+�X���u<1���101W�הּ�2N�A�e�30A#0���"�4N�;2e�5��|�p���"��CalxN �0�O��Z��0�O�$�S�%j{�u��� �0S�}���um�p��\bbk96M8�!68�!��b�.eq969�9�%���F0b�� "BB�OX�ۍ�sch�ed����setau~Xk��� ffH )�0�eq)��0��col(�1bx1c��8�li�Љ� aI���W!i�e@m�{rof$TP EB!lTA&@ry|M427��*l!(T\�Q!RecX"H
�qz�?$it%x�?#сk971�!�71�{�F�$parecjo��A��?'�����Xrail�@nage��~@]�j�D2E� [0 (?:H͒V|x@1ipMa��T�3�p�!4�"4��u��3paxrmr "XRM$��3�rf�Ͼß1�1���0�yturbsp�'G#��^@ �015: ��625t/~A�� \BH�'ZDiy!:k�E�6�"A���H� ��7��P�.�E!pd? "TSPD�}�T�GtsglD��kY`��O�CiCsRct%���HvrvQ���K��P,��A  1q#-a21�Y@AAVM �r�-b0 �fdE`T�UP him (�J545 ly) �i`616 V2VCAM .CLIO Y1�0k 5W` (=F�`MSC ���b�Ps�STYL��Sua28 kr�`N�RE I��`SCH�gRpDCSU� tpsh �ORSR �ua0�4�EIOC�W`\fx�`542� LEX"�`ES�ET��iay`0sh�i`7y`"RMA�SK�b7o�-`OKCO[�x�a7p3Sv( q`t7p0kv6U`xvs39_v�xLCHRvoOPLG�w03;uOMHCR3MpC�`hYaP`�p6�.fia�54; #�MpDSW�`588�ip1�a�37 88 (D�r0c�5r4���r7 qj5r5�5r^v��p5�"9PR�ST VRFR�DMC�S�a��-`9�30 ��`NBA�  g1�`HLB �3 (�aSM�� �Con�`SPVC� Lia20�#-`T�CP aram\TMIL r��PACC�TPT�X �p�`TELON 96�0�r9/u�UECK�1r�`U?FRM etL�a�OR ���`IPL^KeCSXC�pj�q�CVVF l F�7�HTTP st�rbZ0zcpCGy�8~�AIGUI�p�7 ��PGS To�ol�`H863 �dj��qM�Oq3^
vJ684c�\$�@��sق�s'�1ے�s�a96 TFA�Dȑ651�Cq5[3 � oo�b1��44r-�k�r9�V�AT��J775 ��R�6uAWSM|ے�`CTOP ��q�`old��a806;!diy�XYY��0 e��i`885	 '��`L�`u"�`�u 7H�`LCMKP<��pTSS J%��
�W�CPE \�dis�`FVRC� m��NL�U0�02 
�en%�6� 65Jr'�7[�U�0�po�ࠠK���tL� I�4 URI�5��&�U022 ns�e�{�3 APF)I�`{�4�2�`-����alOP��1C�3y3O�͐tptsD`oU040g�43��ٲ4�۰j� "s!w%�1`b	�4�C	�k5 ��wx�57�eOU061��S�6ұrob9�5g�i��C68����!!��7��w�7�Ё�%���"r�key��3w��4�?ǽ���T���8'�0;89�U09���P���9:���2 &�l* �9&�l��9B�Vr�U15�P�M� sl�A �3#�}���1�q�0v4�7��10K8 	�eэphc ���s�1�q�4+�1�����A�5/�tx�1����1]pu�Qѡ�Bt�1�����`��3��
��6��1!p �`��- W8�147? ase C�U`�sB�1 82��1��4�8 (Wa�i��59 ��aU�166�W�1�W�4H� j U�6�#U�7�3�U�8�3ѱ��B��1<{��2 act���?6 "MCR@�ِ�4�1������96=7ǑU193�3��E6��2Y�sP��2A��21��as�F����<�2-���E�2 wF���55�(���U ��cر5)�w�� �q��p����qf��L���$������q4d��2g�8q��8�51�""]� }�q��< b������B]�� f�; �`�̑ � 8 16 (ݰ�BA��A AҰ�]���g :��!��`8 bbf�o=� t� j�� 7 �\� ]��� �2 k_kv��74 &!����W0�H5��57&�5�79 h� L82� %"��4 %3��5����5��<1��594 U21'9 7,-�6�p�Ž6i�\tchH6�ur% �4S3� �90� h�&�\Oj670��q� ��r!tD�4��&ڝt�sg�lc$�S�FrE�H��`#F�����hk$ �� sC�� ��"F�L��dflr0��� �� ����fu!l%�gvPva����sA�����"D��3��!creex���!�%�!�%��,���6j6�s�!prs.�!�%�!�5�hA�P 5�f�sgn��/�/�,at<D�AD���qs`>R svsch`@Q!Servo S�!�uleoCA5SVS�!44���F��1� (�0Ached��0,1�EA၍�� �2Q��0��^�r0�U�)1BBc��� %P5�)Q1�V-#�3�1css "ACS� WVY88"gA�`8!�/�0��@e�Ҿ#M��C�3~�torchm�0n�- TQMa�1x�1M%'�9 J5lA�598 א1�!7)P8<P(1̢A�ء8%R1Qte,�!)E� A5E`ASv�� m�LC6ARC_� 51�4q� �V�Ht!tc�A耥Q�4���R F1 7T!2�SEPBPQf�-!�RtmkQ!p@610X��/�PRC8S�Q�#�S�) P�2a96`xAn`X�D.<bH5�1@�U�}E� T�Qf#`  aQ!<���F!�T!!�aa4�3FcRO�Ttm�R�!av`58�_�WP��M�A$q�E8��>rp�i�n_���o�@e`AcB�rr�)u�!�U�etd�ѧ�U�Qoveto�#$,�S��mmonitr`42�=�Q�c�st,"M_va�P47M��V�0��! 5�q���asmeQ!Ɂrol�Al��43$Q0  S�p��1�01$P25��AKR  �� �0S�(V��Ɂ)xj818\n�l`mD��zN��r�M�PTP"�O��qmocol�]/
�Y1��4Xa�@��2�0i�5�3(1��Touch¤!sؠ�2%qD2J5  !IU�٠��= b�0n��A��]�vP���0z�EOWJ�th���Kwc���{�ett=h8!THSRXâm��t�o "PG�IOsRd�'z�wk�� "WK1�aL&M]H�PH54�5�Q�5�o��m`A��q@7z@6���18�a�PMo\r��tsn�@T�A �o�c���"�����m�uA��T��p���T?�|�m4�T	M�!2�54�>�����m9�w�f��S�3G��qor�3���"64 1���8ⱐQ!A�,HE!pRU <�m��Re�h-g "SV�GN_��(copy "COTA��U(��|r#j0 "FSG���_�eh��f�@w�A�SWwjRbY=sgatu���!�;B�;tp�ATPD7��9 a79s����ssg8!��GAT&o�<Rc9   �Ħ�1�t2`%1�&��1�bpv�1��&��1��B �1� 6�1�c�hr��1�|v�1�s�m��1�v���gtdmenps1�(v0!|1��mkpdt�r`1��]A1��pd���1�$&�1��mvbkup.1��6�A<��mkun��G�spr���mkl1�4e�P�s1�ni��0&�1�ldvr���glg�t�1��&���n#�auth�.p��&��1�����) sud�1�7� 1�G�d1��\1�g b2��p�w 1�6O�Ł4� 1�Ђ   946"1�����1�t\paic\?p4k9471��wc��1�icta�s-�Mpa�c�ck0m	�	g�en!1� wl䟰Q� stfq��q�wb����p�����vri/ �4�^��B1�D���Pflow�@��A�c0ow�3<R5�0?���Q�TR�  (A0e T�)B�Ԗ�cud!�w�1��z�3ac�$046 a� =�f�+paRa���!1�355Ţ1�F��ѡ�)a%��;:af'cald� �&�0P����%�f�m:@�"�#�4�`��'a`"��3U���$�B1�! track���@a�ine/Rail� TrP��{(69�/�@ (L !iEYB �ʔ_VB!Bu���a YB38P�48 '7�	�F2��4��/(�C�B1�3Ţ3�/�fIUal��1�NT��0��VA��zQin�p�?0HVaen0�?DX�WApuA�YqBzQtstd�0U�@1GW  ��]�j�VD���E&���VH@���opene�rs^CO�`�ADev/w'~6�F8���`�����bA�aes�# 1�]�ג�d���하m�d1�k9�@7�6¾�#1��/b�epa;op`aOPN�Wj8�`��Krcel}?�Exg���Y`5Dv��tscx?t��a�s= Fuvrop /�Dw�nDh��bAr5���QB�g�dk�j!�� Pumpv$Aᛑ�@/�1�a;��M�� T�q�i���t4U<�1� 0S��O� \mhplugB�gr7Gh���u|b,Z#��ioh#C{p��\v(�ALIO1�1�@M7��93�Q51��91�����4�� S�T�
R�t�J9899��/RLSE�g1ʖ@Cd�(M�1�/O��'�Q�)�D��G1 0zq�H155'?��|zq�tcmio���MIO�$�tc>�q"CL01�UQYcP�|�io��u~0%�l9�zp��v�"1o���Q�tzt����dtz5I$��V%<�rh#Inte�Q��� Co~Po�qvR�P1�hd�B554 (l�oBv�,�Q�H���Tcipc�oo�ڱp	5�A�(
�������D�"7`���aڰd�QCD�W�	����p8��ڱ�rcnd�_׳1p�a�ײ� �����S��a��OƳ2kz�rpcCrt�ᱯ�pٱdEc ��S d�\���u�E!<߳vr2k�pE �A�-�x�_B\"� choO�l"uC��Y 1���630@ᗷ�@��� �ӿ�q��ԑ�GT�X�? �Е1chpC "��XOh:�3��&�"5x!E��\p3� ���P��j�d 1`1�$h��Plo���ұ�ch��3���s1��a�01 ���#Ar��0� !oCB��spq[Jm:�k�7�)�vr�Ҿ���a!X%�-J�FRAJ�Watpqrnev'������fQ��D5�`��KrboT ,�$���PG�[!�sm�ICSP\QQP5y�<�!QP���nj�H51z�93QP	7y�6��������5��R6QP���N�PR�`(P@aam S`u�b��ĉa4tpprg�p�B�	��Z�qratk93�2(q v��sc� "iC��~�atpr�_�qqz�;F��LGdsblfl�t{�ёsableO Fau`��CPa�v�aQ��`aDSB' (Dt$�t�d�A ����QPh"�E1��`f$�*��3[S� A�"tdj  "PaV�Ohf$��1sbj!��1�"\�:1gc��.�f%�du�5�50^CAdjust Point�b��J/��-�0�4�a�昐A��j�O�N0\�sg�4��w�1\�ada��"ADJ��M�j0�etsh=am�SHAP0���XDjpo �e��G�a���UGQPG'.��1:�kr@ab5�J�KAR`��iagnosti���!�a��66 JP�C��a=P(QL�Q�&T�o�fkrlde P@���	 ��SQ���)�3/ρ[pp��D'BG2t�!O �U�R ѯ#��V��F( �шSX7��Q�ip{�M��ipper Op�Pq����78 (MH Gw�1Rlbk_ �fTcBQ��0&�d038<B8t��E��c
�9_9t��Tc��	k����8$q�Sdr npVǁ��Qd�Ő6�Tea�=���r Mat.Handlv ��an`W�� MPL!Gv�A_�p�q(�sє �f����g��b�� a���f������>@ $w����Dw��EI d����uu�m���f�hnd "F�� � ������#� ��p��>��(Pa�0To@�$V�!!�
3#p��a>��{�Q�/k925��26�q�$3�{�p����2	ş��y���gse>0GS �qďėPR��T���a���tp����{�dmon_�q�Ŗ�a3ns���vr��{߀=�����ͪ�<y��wsul� � pen���D��Y�WA��823X�Q
�G�0!'�&P���8QqIQ�GQ �\sl��!q��v� ���������֐�_�`|����"SEDGiO�ٳaQ�tdg�@T �AF8�F���BN���À�Qm�7���ڱA��g�;Ж�Q�����q�S�ileg�y�e���ϟ��9�F'QQ�LaQQj5C17So�3-[JV� ?�'�#4A�49G�A�WL�aw {�no0�Qfԫo�H17D��#a�����0t� � >���LANG j�A�5��5�5� ga�d5��C5�TC5�jp� .5�ce���5�i�b=�5��#5���pa�5��C5�WҸ�j53g9.f5�]QRu5�? Env
5�5S���K�3y ��J9 $5�.� �;��G
5�2D25�JS��p�(K}�n-Tim ��"���"��3H�ܹ���\kl5�UT�IL"�����r "QMG��,q5�C5��1 "5�ړ5�|�s5�\kcmn��`+��r5���utM�>_�lread���Cex����"��\��l$"��135�rt[! -5�tuva��л`_��5� �`CV����\p ���Bzp9tbox��<_qcycs}k�RBTvveri?OPTNv��l��e��K����hg/�agp�.v1$�"1$ptl�itDPND��BPm$dn#te\�cym$8$o"��#m�nu3�/�/�/�.5��/�/m$��UPD�T ite��.3 �swto95]�-4oolBD5wb95��-4`FR-4Y�� /2grd�@-4��-4�b-4��w-4 B-4.3��-4�-4 '�-4�.3B0l� /2bx "�5�Q5I.3tl�7��AE�#/2r l\�6�@O�-4\ :4ColD5eMa-4+�C�5K�-4W�Q5�ml�-4Chang�95}�95�qQ5rcm dE�b�OZ�`6�5,r�7�6��7�5&r_+]22=_O]2� c_u_23U4<_N^57�_�_1UCCFM�Ey��_accdau59#�6cAEX`�/2|�Da��4|aO/Jm�a�5� -4@�4�aAOSJ	Q�e �o�oY��-4��ZDQ-4sk��?�@rtet�q-4\$�3�q�eunc.-4��4�q�5sub�5��5E�q�5cce�@oRf@^opm4E�o�fv�7 �o�eT �c�o�nt$
Pte;�q �@�f\���k��6;�-4Ѓ -4K�D��zh!-4xmov�b�q��et���f�"�tg?eobdt.������etu� ɐ��ɐ���tɐٓxߟ�z���var'��x�y&��pclJ�c�ɐ��ɐ�eɐgr�ipsu����ut�i�����infp!o��ܯ�ɐ������\����ɐ�Ʊ�
8�p��n��ɐ%�ɐZ�mT���ɐԶ��\�ogġ�Ʊ�%�p�\�Gpalp�����s�����ɐݵ��Ŵ����px�p����pkagd�|%�7�lclayY�k�A�ɐ��dɐ5�p�������B��|�|�Ⱥ�����q����rd9mͿ��rinT�-߂?�sO�Q�c�̿޼s����ߧ�tv�ߧ�h8���stn[`�J�tX01ɐ)�Dɐ� �Tul4�q��rg�26Ϥ�upd�����vr����נ1�}�3�נ��ϵ�il3C�U�l4����T�5e�w�s ߘ�֠�ߎ��wcm�(��x�ferϪ�tlk�2pp��con9v�朗cnvݑ���5�ag, y�lc�t���n�p��nit0���d���(���  �ɐ 0S�(V�U69al �pm�Wse��2����V� C��(�z���A�0�|�m����&$��޷'#ro��T/f(&���p1�mI��,��$� �+���/�)G�?�+ �� �L�ɰm ∡ P?b6D�4rg�� ���������?�9��  O�7������ >�/�T�a�8/�C�� ���E��b,֡)?�*��nq?_9l�-!H���  �HA �|�p�QU1 �p! O���P ���S 	�Q�R@�t�`  ?���ɐ8� �M�.O�reg.ԃnO�o�99 �� ����$FEAT�_INDEX  ��S ����P�5`ILEC�OMP >�{��baPa��RUcSETUP2� ?belb��  N �aUc_�AP2BCK 1�@bi  �)8�R�o�o  %�o�o�Pe`�o)oe�oU �oy��>�b �	��-��Q�c�� �������L��p�� ���;�ʏ_���� $���H�ݟ�~���� 7�I�؟m����� ��� ǯV��z��!���E� ԯi�{�
���.�ÿտ d�����Ϭ�*�S�� w�ϛϭ�<���`��� ߖ�+ߺ�O�a��υ� ߩ�8߶���n��� '�9���]��߁��"� ��F�����|����5� ��B�k��������� T���x���C�� gy�,�P���qi�`P�o 2>�`*.VR�H� *Kq�w���2PC��� OFR6:���/�T@`@/R/�=/�|,C`/�/�*.F5�/�	��/ <��/$?�+STM @D2M?X.�E?�=� �iPendant Panel�?�+Hz?�?j7�?�??-O�*GIF7OaOl5�MO
OO�O�*JPG �O�Ol5�O�O�O5_��
ARGNAME�.DT?_�o0\�S__� �T�_@_	?PANEL1�_�_%o0�_o�?�?�_2orog`oo/o�o�Z3�o�og�o�o�oH�Z4zgh%�7�KUTPEIN�S.XML�o_:�\���qCust�om Toolb�ar(��PAS�SWORD���FRS:\k�*� �%Passwo�rd Config��������+�� O�ޏs������8�͟ ߟn����'���ȟ]� 쟁��z���F�ۯj� �����5�įY�k��� �����B�T��x�� ���C�ҿg����ϝ� ,���P����φ�ߪ� ?�����u�ߙ�(ߒ� ��^��߂��)��M� ��q����6���Z� l����%����[��� ������D���h��� ��3��W����� �@��v� /A�e���* �N�r�/�=/ �6/s//�/&/�/�/ \/�/�/?'?�/K?�/ o?�/?�?4?�?X?�? �?�?#O�?GOYO�?}O O�O�OBO�OfO�O�O �O1_�OU_�ON_�__ �_>_�_�_t_	o�_-o ?o�_co�_�oo(o�o Lo�opo�o�o;�o _q �$��Z �~���I��m� �f���2�ǏV���� ��!���E�W��{�
� ��.�@�՟d������ /���S��w�������<�ѯ�Ơ�$FI�LE_DGBCK� 1@��ʠ��� (� �)
SUMM?ARY.DG篓�OMD:�[����Diag Su�mmary\�i�
CONSLOGQ��4�F���߿n�Co�nsole lo�g�h�G�MEMCHECKտ��J��c��Memor?y Datad�l�ߑ {)O�HADOWY�>�P���t��Shadow Changes���£-��)	F�TPҿ?���C�n����mment T�BDl�l�0<�)�ETHERNE�Taߑ�"�����n��Ethernet� ��figura�tion��s�V�DCSVRF`�F�X��q�t�%6� v�erify alylt�£1p�1�DIFFi�O�a����u�%��dif!f���"�6�1������{� �����{	9�CHGDE�W�i���u��&���9�2������� 1�����GDM_�qu�.9F�Y3���� 1���GDUg�y/u�6/��UPDATES.�U ;/��FRS:�\S/�-o�Upd�ates Lis�t�/��PSRBW�LD.CM�/���"�/�/��PS_R?OBOWEL��g� \?n?���?���?�?W? �?{?O�?	OFO�?jO �?{O�O/O�OSO�O�O �O_�OB_T_�Ox__ �_+_�_�_a_�_�_o ,o�_Po�_to�oo�o 9o�o�ooo�o(�o !^�o���G �k ���6��Z� l�������C���� y�����D�ӏh��� ����-�Q������ ���@�ϟ9�v���� )���Я_������*� ��N�ݯr������7� ̿[�ſϑ�&ϵ�7� \�뿀�Ϥ϶�E��� i���ߟ�4���X��� Qߎ�߲�A�����w� ��0�B���f��ߊ� ��+���O���s���� ��>���O�t�������$FILE_ {PR� ����������MDONLY 1�@���� 
 �5�Y�0}�=f /����O�s �>�bt �'�K���/ �:/L/�p/��/�/ 5/�/Y/�/ ?�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO��O
_��VISBC�K������*.V�D_[_�@FR:�\F_�^�@Vi�sion VD file�_�O�_�_ �Oo�O)o�_:o_o�_ �oo�o�oHo�olo �o�o7�o[m(�  �D��z�� 3�E��i�����.� ÏR���������A� ЏR�w����*���џ `����������O����MR_GRP 1�A��L4�C4�  B�9�	 ��񝯯����*u����RHB� ��2 ���� ��� ��� ݥ���������ި%��ߤA�5���_�J�K�t7I�TWH�h��T���R��*P��M����q� F�U<�Hp�G,*�;��h;r���@N�-��@�������E��� F@ %5�U1ŝ�J��NJ�k�H9�H�u��F!��IP�s��?@�u�ÿ�9�<9��896C'�6<,6\b� ������������ ��A9�A�?�M��r��ߖ߁ߺߥ�  >�o"A\a@��@���� �����8�#�\�G�� k���������4�;BH9� ��8������>�P�`�
��P�X�P�k(`�w�����B�����M�O@�33������\��UUU!U<��	>u.�?!���k�����=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!��7�:�7p��D��@ D�� CY�@�UC���Ώ�'�������-�/ �C/�#/1��/Y�/ �/�/�/�/�/�/0?? T???x?c?�?�?�?�? �?�?�?OO>O)ObO MO;�N�P�^O�OZO�O �O_�O+__(_a_L_ �_p_�_�_�_�_�_o �_'ooKoXi�Xo~o �o�oi��o�o=o�o�o BT;xc� �������� >�)�b�M���q����� ����ˏ���7�/ {/%/7/��[/��/ܟ �� ��$��H�3�X� ~�i�����Ư���կ ����D�/�h�S��� w������O㿩�
ϥ� .��R�=�v�a�sϬ� ���ϻ�������(� N�9�r�]ߖ�]o���� ���߷o�{�$�J�5� n�U��y������� �����4��D�j�U� ��y������������� ��0T�-��Q� �u������ϟ5 GP;t_��� ����//:/%/ ^/I/�/m//�/�/�/ �/ ?ǿ!?�?Z?E? ~?i?�?�?�?�?�?�? �? OODO/OhOSO�O wO�O�O�O�O��
__ ._@_�d_�O�_s_�_ �_�_�_�_o�_o<o 'o`oKo�ooo�o�o�o �o�o�o&J5 nYk�k}�� ���1��U�� ��y���ď���ӏ� ��0��@�f�Q���u� ����ҟ������,� �P�?q�;?��[��� ί���ݯ��:�%� ^�I�[��������ܿ ǿ ���6��OZ�l� ~�E_Oϴ�������� ���2��V�A�z�e� w߰ߛ��߿������ �,�R�=�v�a��� ��������'�I� K��7�9�?���o��� ��������8#\ G�k����� ��"F1jU g�g������/ �/B/-/f/Q/�/u/ �/�/�/�/�/?�/,? ?P?;?t?�?MϪ?�? �?���?Ok?(OOLO 3O\O�OiO�O�O�O�O �O�O�O$__H_3_l_ W_�_{_�_�_�_�_�_ o�_2oDo�eo/��� �oe��o���o��
%o .R=vas� �������(� N�9�r�]��������� ޏɏ��׏8�ӏ\� G���k�������ڟş ���"��F�1�C�|� g�����į�?ԯ��� ��?B���;�x�c��� ����ҿ������� >�)�b�M�_Ϙσϼ� ����������:�%� ^�I߂�Io[o��o�� �o�o��o3��oZ�u� ~�i���������� �� ��D�/�h�S��� w�����������
�� .����'�s� �����* N9r]���� ���/ۯ8/J/\/ n/5��/��/�/�/�/ �/?�/ ?F?1?j?U? �?y?�?�?�?�?�?O �?0OOTO?OxOcO�O�O�O�O���$FN�O �����A�
�F0Q P T�1� D|���@RM�_CHKTYP � �@����@���@�QOMP_�MIN"P�����NP�  X�@S�SB_CFG �B�E ��{_��rS�_�_�E�TP_DEF_O/W  ��-R�X�IRCOM!P�_��$GENOVRD7_DOCV���l�THRCV ded�d_ENB�_ �`RAVC_GR�P 1CdW�Q X�O�o�O�o�o�o�o �o&J1nU g������� "�	�F�X�?�|�c��� ����֏������0�.bROUp`I�HQP�����R��8�?T쀟3��|�������  Daڟl���@@�B������o�4�g`WSMTmcJtm�𗯩����AHOST�C]R1KO�pP�Ya� M������0�  2�7.0G�10�  e'�t��������� b�ۿ����4�˿ų�	anonymous8�f�xϊϜϨ����л���%�'�� [�0�B�T�f�x�ǿ�� �������Ϗ�E��,� >�P�b���������� �������(�:��� ^�p������������ �� $s���� ��������� K� 2DVh��� ������5GY km7/�v/�/�/�/ �/�/�/??*?M/ ��r?�?�?�?�	/ /-/OA?c/8OJO\O nO�O�/�O�O�O�O�O OM?_?4_F_X_j_�? _�?�?�__%O�_o o0oBo�Ofoxo�o�o �o�__!_�o, >�_�_�_��o��_ ����So(�:�L� ^�p����o��ʏ܏�� �u�١ENT {1LO� P!��.E�  A�3�p� _���W���{�ܟ��� ß�6���Z��~�A� ��e�Ư�������� � �D��h�+�=���a� ¿��濩�
�Ϳ�@� /�d�'ψ�KϬ�oϸ� �������*���N�� r�5ߖ�Y�k��ߏ���������QUIC�C0!����p�3�1 q�M�_���3�2�������!ROUT�ER�����`�!�PCJOGa�<��!192.16?8.0.10:��NAME !"�!ROBOT����S_CFG 1�K"� ��Auto-st�arted`tFTPkH���s ������$� '9\J��� ���Jv!3E/ Y{1/b/t/�/�/g �/�/�/�/?'/�/:? L?^?p?�?�?Qcu �?? OO/$O6OHOZO )?~O�O�O�O�O�?kO �O_ _2_D_V_�?�? �?�_�O�_O�_�_
o o�O�_Rodovo�o�_ �o?o�o�o�og_ y_�_1�o��_�� ����o�&�8�J� mn��������ȏڏ );M_a�F��j� |���������֟��� �/�ɟßT�f�x��� ������!�#��W� ,�>�P�b�t�C����� ��ο�����(�:� L�^ϭ���ѯ���� ��� ��$�6��Z� l�~ߐߢ���G��������� ���T_ER�R M��.�>�P�DUSIZ  j �^���U�>n�?WRD ?����  guest\��������������SCDMNGRP 2NwX�����p��\�KM� 	�P01.14 8~��   y���}�B   � ;���� ������������������?�����~��\�������|����  i  ��  
���ҕ������+�������
���l��.؋�"��luop 
dy�����|��&�_GROU8�]OM� �	0��p�07�	QUPD'  ��U��!�TY�M�@�T�TP_AUTH �1PM� <!iPendan������!K?AREL:*���KC�����VISION �SET� ://�� �Q/?/i/��/{/�/ �/�/�/�/"?�/>YCTRL QM��P�v5��
��F�FF9E3.?���FRS:DEFA�ULT�<FA�NUC Web �Server�:
 Y���A<OO*O<O�NO`O<�WR_CONFIG R<�� �?>�IDL_CPU_PC�0���Bȩ��@�BH�EMIN�L���D?GNR_IOG�|����S�@NPT_S_IM_DOV[�TPMODNTO�LV 3]_PRT�Y)X�B�DOLNK 1SM����_�_��_�_�_�_o|RMA�STEP&|R_O�_CFG"o4iUO�DEo6bCYCLE�do4d�0_ASG s1T<���
 o �o�o�o�o!3E Wi{���k�bNUM{�Q��08`�IPCH�o58`R?TRY_CN�0
R<Q�6bSCRN>{㊗Q�U� 6ba`?b�UM��p����$J�23_DSP_E�N� M�ᆀOB�PROC��LUMiJ[OG�1V�@Q�?8�?��{���?ŃPOSRE���VKANJI_@`d�
_H��V�W�L�}6h�1�C�CL_�L�@�r�H�EYL_OGGINB`����Q�PLANGU�AGE �6�Be�4 �>�LGW�YXf?�ҧ���x% ����?��@���'�0��`$�>M�C:\RSCH\�00\�?�N_D?ISP YM��p��|�z�<�LOCGR��BDz�DA�OGBOOK Z�k�R�P�T�X ��B�T�f�x�������1����v6	�<��⸥���_BU_FF 1[�]� I�2��H�S�h�d�n� �ϒϿ϶��������� +�"�4�a�X�j�|ߎ���߲����ߔ�ˀDC�S ]� =��;���C��5Y�k��}���IO 1^��k t��� � ��������� �2�D� X�h�z����������� ����
0@Rd�x��EPTM  GdR2���� 0BTfx�� �����//,/8>/)Ĩ SEV:���]�TYP��`�/�/�/ �-�RS�0���*�2�FL 1_��@��9�9?K?]?`o?�?�?�?�/TPѐ��"ݭNGN�AM��p�tU�UP�S��GI���E��A_LOAD��G� %��%��_�MOV[�aO�DMA?XUALRM�w�@�x{@AdQ:�<��C��y@C��`��Oj��lM�@̀Ҁa�k ��X�	�!�p+e���OΤ,RX_C_U_ �_7�|_�_�_�_�_�_ oo;o&o_oqoTo�o �o�o�o�o�o�o�o 7I,mX�t� �����!��E� 0�i�L�^�����Ï�� ���܏��A�$�6� w�b�������џ���� ������O�:�s�^� ������ͯ���ԯ� '��K�6�o���d������ɿ�GD_LDX�DISA�0���M�EMO_AP�0E� ?a+
  � ѹ%�7�I�[�m����ϣ�y@ISC 1ba+ �����'T ,���
ߺ�C�.�g�N� �ߝ�߬߀�����	� ��?���N�"��� ������b������ ;�&�_�F�������� x�������7�� F�|��� Z���3W> {��p����/��_MSTR �ca-%SCD 1d͠�m/��/ |/�/�/�/�/�/?�/ 3??W?B?{?f?�?�? �?�?�?�?�?OOAO ,O>OwObO�O�O�O�O �O�O�O__=_(_a_ L_�_p_�_�_�_�_�_ o�_'ooKo6o[o�o lo�o�o�o�o�o�o �oG2kV�z �������1���U�@�y�/MKC_FG e--��~<"LTARM_���f��� �v������METsPU�n���5)�NDSP_CMN�T�����#�&  	g-.a�v���y����#�POSCF/��:�PRPM.� �PSTOL 1h��{4@��<#�
�� t���������/� q�S�e�������ݯ�� ѯ����I�+�=���i�#�SING_C�HK  ǟ$M/ODAQӃi��a������DEV 	�K*	MC:�HOSIZE�--ȹ�TASK %K*�%$123456�789 V�hŷ�T�RIG 1jK+� lK%%�a��� � ������M#8�YP�#���5$��EM_�INF 1kڇ� `)�AT&FV0E0���a�)I�E0V�1&A3&B1&�D2&S0&C1�S0=P�)ATZaߵߜ�H����p���	��A�9���]�D��� G߸�k�}� �ߡ����6�m�Z�l� ��K����������� �� ������hs�-� ����}���� @Rv);M _���+/*/� N/	/r/�/k/�/[m �/���&?8?�\? �/�?;?E/�?q?�?�? �?O�/4O�/�/?? �OA?�O�O�?�O�?_��O_B_)_f_��ON�ITORJ�G ?���   	EOXEC1p��R2�X3�X4�X5�Xy��VU7�X8�X9p��R 0Bd�Rd�Rd�Rd �Rd�Rd�Rd�RdPbdbc2h2'hU23h2?h2Kh2WhU2ch2oh2{h2�h�3h3'h3�R��R�_GRP_SV �1��>ї�(q�������Yp�?��=
҅?�?OȽ�f��@��_DR&Λ�PL_NAME !���p�!Def�ault Per�sonality� (from FwD) ��RR2-q� 1m)deX)�dh��q7�X d v� ��$�6�H�Z�l� ~�������Ə؏����� �2�D�V�h�t�2 �������Ο�����(�:���<��d�v� ��������Я������*��R,r 1r�yհ\��, ������f� @D7�  z�?���f��?������A'�6xz�ܿ��;�	l���	 �x7J԰������˰ �< ���� ��IpK��K ��K�=*�J���J?���JV尻�"�ɱT��:�L�Ip�@j�@T;fb��f�n���%�4���=�N�����I��g��a������*��* � ´  ��PÕ>�������n�?z���n�Ͽ�Jm����  
�ғ�%��Ī�9���� �`�  �P}pQ}p�}p| � �r�/׈�+�	�'� � ���I� �  {��J�:�È��?È=�����6����	�ВI  �n @
�+�l�$��l���9�A�7�yN�p|�  '���_���@2��@�ӹ�f£�@��C���C�pC�@ C���C��C��o�
��A�q��P� @���
0�B�p*�A��2���a`�o�R�n�Dz�ˀq��߁�������2���( �� -����������No� ���!�o��M� �?�ff ���/A�� ��v�7�a��
�>��  P��2�( o��e�����ڳڴ^D�?��o�x"�Ip<
6b<���;܍�<����<� <�&�KNA둳��|nO�?fff?��?&�3�@�.���J<?�` �M����.ɂ�� ���lƴa2//V/ A/z/e/�/�/�/�/�/�/8�F�p�/4? �/X?�y?�K?�?�ȿE�� E��G+� F���?�? �?O'OOKO6OoO.�BL��B�_0��� �OUO[��OcO_o?5_ �?\_�O�_�_�_�_U
��h��V�W>��r_on_/oo,o�eo�GA��d;���C�Ro�oNoD����ؠ�o�o%5yķD���8C|�spCH�5"Z�d����a�q@�I�~N'�3A��A�AR1A�O�^?�$�?���;��±
=�ç>����3�W
=�#��n�{e��n�@������{����<���~(�B��u��=B�0�������	��H�F�G����G��H��U`E���C��+���I#��I��HD��F��E��R�C�j=z�
�I��@H�!�H�( E<YD09ڏ�׏� ��4��X�C�|�g�y� ����֟������	� B�T�?�x�c������� ���ϯ���>�)� b�M���q�������� ˿��(��L�7�I� ��mϦϑ��ϵ����� �$��H�3�l�Wߐ� {ߴߟ߱�������� 2��V�A�z��w�� ������������tR��q(�q���������e���v����a3�8�x�����a4Mgs�������IB+���a���{�& &	fT�x���e%P�P��A�O	�\���*<��R�^p�����  ����*//N/ </r/�)�O� ��/�/�%�Q�/�/�/?8?'?9?  N?l/��?�?�?�?�?�2 �F�$�Gb����A��@a�`rqC��C@�oTO� q�{O�F� Dz@��� F�P D�!�]O�O�I�cO�O��O__1_�c?��W�@@8Z^4� �� �� �n
 8_�_�_�_�_�_ �_oo+o=oOoaoso��o�zuQ ������1��$MSK�CFMAP  �R5� �`6uQqQ�n�cONR�EL  ���a� �bEXCFE�NBw
�c�e qF�NC'tJOGO/VLIMwdpr]d�bKEYwsu]�bRUNc|su��bSFSPDT�Y�p)vu�cSIG�NtT1MOT�eq�b_CE_�GRP 1sR5�c\:�I�2�m�� �Di���a�Ώ��Ï� ��(�ߏ�^������ K���o�ܟ��ɟ �H���l�~�e���Y��Ưد�����F�`TC�OM_CFG 1�t�m�V8�J�\�
��_ARC_$r��2yUAP_CP�L��6tNOCHE�CK ?�k �׸տ���� �/�A�S�e�wωϛ��Ͽ������kNO_?WAIT_L�w�e6�NT �u�kw[�5�_ERR!�29v�i�� ��߲߾��c���ߴ��T_MOc�wj�,� '��3���P�ARAMd�x�k�tV#���=?��� =@345678901�������� ����+�U�g�C�����y�������t����UM_RSP�ACE�olV>H�$ODRDSP���v2xOFFSET�_CART��yD�IS�yPEN_FILE� jq^�+��v�OPTION_�IO�YPWOR�K y'�5s x�fRuQ��2��2	 �	2���[ RG_DS�BL  R5s�x\�zRIENTkTOp!C�oP��a.A[ UT_SIM_D��b�b[ �V_ LCT z�?�*+^�)�_P�EXE�,&RAT�8 jv2u�p0"� UP� {.�PS0�`�/�/�/�/�)�$O��2 �m)deX)�dh��X d��?-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�H2
?�O�O�O�O�O_ _1_C_U_%�<�O_ �_�_�_�_�_�_�_o@!o3oEo�O� �Ov �1r(���(���07�, �lp�` @D7�  �a?��c�a1?m�a%�D�c�a����l;�	l�b	� �xJ�`�o�u��`� �< ��	p� �r��H(���H3k7HS�M5G�22G�?��Gp
��������Yk|��CR�>��qȋs�a�����*  ���4�p�p��pT����B_���{�j%��t�q� )�/��aD�������6  ����P� Q� �� |�Б�������	'�� � ͂I�� �  �=�i�=��������a	���I  ?�n @)��mC���m��[��9N���  '� ��t~q�pC�C�@�s��pC���ҟ 5�
S��=x@#�7~�9�^�n�B�I�A8��Q��� 0�q��bz比������ȯ�����( �� -݂*�΁06���Am� �0rx���m�lp �?��ffU ܫN�`����n�8m྿̺�>�  P�aզ( m������� q�c�d^#?��m�xA��n�<
6b<���;܍�<����<� <�&1j�m�A0��c�|��n�?fff?0��?&����@�.��J<?�` ��l�����dѩ�e�� �gߋ��d��Q�<�u� `ߙ߄߽ߨ������� �)� �M�8�q���
���j���f�E�� �E�0�G+� F������� �F�1�@j�U���y�[bB��A��|����t�z� ��3��T��{������t��h��<u�w�>��*��N9K���A��Z�_�Cq�mc��?��//D///T)���pٞ�aF�`CHT/A
$� �!�!@Iܝ�'��3A�A�AR�1AO�^?��$�?��������
=ç>�����3�W
=�s#�>��+e�� �������{�����<��.(��B�u���=B0�������	3�\*H�F��G���G���H�U`E����C�+�Y-I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0X/�?O �?/OOSO>OwObO�O �O�O�O�O�O�O__ =_(_a_s_^_�_�_�_ �_�_�_o�_ o9o$o ]oHo�olo�o�o�o�o �o�o�o#G2k Vh������ ��1�C�.�g�R��� v�����ӏ��Џ	�� -��Q�<�u�`����� ��ϟ���ޟ��;��&�8�q�\�(��ٙ�,�����]��������p!3��8���ӯp!4Mgqs����IB+��+��a���{�E�E���s�����Ϳ����Pe�P�� (�{�4��I�[�իR}Ϗ��ϳ�������  ���˿I� 7�m�[ߑ��H� ߿������������"�4�F�X�   m�ߵ��������缿2 F�$�Gb��ϲ����!C���@�s������ F� Dz�/�� F�P �D�����������,>P�?_���@@W
}����������
 W��� �&8J\n�����*� ����˨�1��$P�ARAM_MEN�U ?q���  �DEFPULSE��	WAITT�MOUT+RC�V/ SHE�LL_WRK.$�CUR_STYLv G,OPT]�N]/PTBr/l"CB/R_DECSN  ��,�/�/�/
??? )?R?M?_?q?�?�?�?��?�?�USE_P�ROG %�%��?#O�3CCR ���6G_HOST7 !�!;DxO�0JT�BO�C[OmA��C�O/K_TIME�"�B�  �GDEBUG�@��3�GINP_FLMSK�O(YT��9_*UWPGAUP \���g[CH6_'XTYPE����?�?�_ oo#o5o^oYoko}o �o�o�o�o�o�o�o 61CU~y�� �����	��-��V�Q�c�u���*UWO�RD ?	{]	�RS��	PNeSW�V$ڂJO�!΂�TE�@�VTR�ACECTL 1�|q�� ��� ����4��DT Q}�q�c�(�D ȿ  L� �p�Mt�� v�O� ��� ��� ��� ������p�Et�t�V�v�t�t���v�t���v�� v�t�t��v�TN�v�!t�"t�#t�T'�v�%t�&t�'t�(t�)t�*t�@�v�U,t�-t�.t�/t�U0t�1t�2t�3t�U4t�5t�6t�7t�U8t�9t�:t�;t�U<t�=t�>t�?t� n v�]�v�� v�� v�Dt�Z v�Ft�Pv�Ht�It�Jt��Pv� s��������Q�������သ� ��U��V���W��X��Y��Z���[��\��]��^���_��`��a��b���c��d��e��f���g��h��i��j���k��l��m��n���o��p��q��r���s��t��u��v*��w��x��y�������&�֘� ;Ҙ�#Ҙ�KҘ��P��P� ��� ������U	��
�������������@��������۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y���l� Е����������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_Е���_o"o4oFo Xojo|o�o�o�o�o�o �o�o0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
���_@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n����� ���������"�4�F� X�j�|����������� ����0BTf x������� ,>Pbt� ������//�(/:/L/^/h!�$P�GTRACELE�N  g!  ���f ��|&_UP ~�����!� �!�� |!_CFG �%�#f!�!���$� �/�/;�"D�EFSPD ���,1�� �| I�N� TRL ���-f 8�%G1PE�_CONFI� �>�%��!�$]<LID�#��-��4GRP 1�܂7�!�g!A ����&fff!A�+33D�� D�]� CÀ A)@6B1�f d�$I�&I�1�0� 	 �?�"�+@O ´yC[ODKB|@�A�OmO�O�O�O�Of!>�T?�
5�O4_F^�0_ =��=#�
K_�_G_�_�_�_ �_�_c_�_&o�_6o\oGo  Dz�c�of 
qo�oao�o�o�o �o0T?xcu������IK
�V7.10bet�a1�$  �A�E/�ӻ��A f ,�?!G�^C�>��+���0�T���+�BQ�c�A\i�T�D;�*{�p�"�B������Ə؏�T�O'O�2�8��\�G��� k�������ڟş��� "��F�1�V�|�g��� ��į���ӯ���	� B�-�f��ov���K��� ���������>�)� b�M�rϘσϼϧ���x���=�F@ � �'�۫%Wك�W߉� �ߑ6��������� %��I�4�m�X��|� �����������3� �W�B�{���x����� ��������S ~�w�8���� ��+O:s ^������
�<� //R�d�v�l/~/�� �/��������/�#? 5? ?Y?D?}?h?�?�? �?�?�?�?�?O
OCO .OgORO�O�O�O�O�O �O�O	_�O-_?_jc_ u_$_�_�_�_�_�_�_ �_oo;o&o_oJo�o no�o�o��(/�o b/P/&Xj�/��/ �/�/�/��o��3� E�0�i�T���x����� Տ��ҏ���/��S� >�w�b�������џ�� �����+�V_O�a�� ��p�����ͯ���ܯ �'��K�6�o�Z��� �o�o�o޿*< nD�rk�}Ϩ�� ��φ������
�C� U�@�y�dߝ߈��߬� ��������?�*�c� N��r�������� �0���;���_�q�\� �������������� ��7"[F���� ο����(�0 ^�Wi�Ϧϸ�v� r��/�///S/ e/P/�/t/�/�/�/�/ �/�/�/+??O?:?s? ^?�?�?�?�?�?�?� O'O�?KO6OoO�OlO �O�O�O�O�O�O_�O _G_2_k_����_ �_�
ooJCo Uo����oL_�o�o �o�o�o?*c u`������ ���;�&�_�J��� n�����ˏݏO�� 7�"�[�F����|� ����ٟğ���!�� �W��_�_�_�����_��_ o���6b�$P�LID_KNOW�_M  bd��j�#�SV� �3e=�:e��z����� 7�¿������j�vmC��M_GRP 1�TP��`d�bd@I�)߶B�_�
�_� ����t��@ǘϾ�^� ���ϮϪ�
�����F� �d�(�Zߠ�^����� �߶����*��� �f� $�L��Z�|������`����,�>�#�MR'�ŉ.�Tg���  㢞������������� ������Q+%7� �������� �M'!3���`����Y�ST'��1 1�3e3 �vi�0:o A >/ g�</N/`/r/�/�/�/ �/�/�/�/?C?&?8? y?\?n?�?�?�?�?�?�	O'2(.:/j��<=O.3'O9OKO]O!#4vO�O�O�O!#A5�O�O�O�O!#6_&_8_J_!#7c_u_�_�_!#8�_�_�_�_!#�MAD  wd�3#x`$PARNU/M  ++�5o�"SCHOj ]e
�gpa�i=��eUPD�po�e�t"_C�MP_$�R`ؠ`'�;�)tER_CHK7u��;�Or4�F{RS|�2�#�_M�OQ`��u_�be__RES_G' �+- O���H�;�l�_� ������Ə���ݏ� ���w&@�|�5� �uu@R�q�v��s�@�� �����sPП����s bP�.�3��s�PN�m��r��s `�������rV� 1�P���b@c�X��p�$@c�W�(��(�@@c�V�4���rTHR_INR|�Tau�d<�MASSI� �Z]�MNH�{�MO�N_QUEUE ��.�bvg��g�*bdN.pUrqN��`{�ΰENDб��EcXE����`BE��|ڿ˳OPTIO׷��{ΰPROGRAoM %��%Ͱ�믖o̲TASK_�IQd@�OCFG �����o����DA�TAe���@�2�N�`�r߄ߒ� <ߵ������ߖ��!��3�E�W�
�INFO
e�"ݘ����� ��������)�;�M� _�q����������������n�z�"� �!���OpDIT ����s�WER�FL��#RGA�DJ �b
AЄ�0�?��P��I�ORITY��av�>�MPDSPX���U����OG$ _TG� K���E�TOE��1�b� (!AFD�E��p��!tc�p��!ud|��?!icm���FXY_����b���)� *0J/\/` ���G/�/ k%w/�/�/�/�/�/? �/2??V?h?O?�?s?��?�?*�PORTT3�Rc���u��_CARTREP��bk@SKSTA����zSSAV����b
	2500H863(�ς5D1U�b`@������s�O�O�G	PURGeE�B�	�yWF�@#DO��$�evW�T��a�:WRUP_DELAY �b>TR_HOT{���%o�_TR_NORMAL{�}_�_�VSEMI�_�_oCa_QSKIP1��u;�Cx 	bO\o \@Jo�o�o�ojh�u�o �g�o�o	�o?- Ou��_��� ����;�)�_�q� ��I�������ݏ�� Ǐ%��I�[�m�3�}������ǟٟ�ͥ�$�RBTIFR�R�CVTM.+D��	�DCR1c�8l��qiC ��>��� >�k��o ��U	��I�i��nro¯���<
6b<���;܍�>u.��?!<�&ǯ���)�ŰHB� T�f�x���������ҿ ������>�)�b� Mφ�qσϼϟ����� 5��(�:�L�^�p߂� �ߦ߸���������� ��6�!�Z�E�~��s� ����	������ �2� D�V�h�z��������� ������
��.R dG������ �*<N`r �o�����/ �&/	//\/��/�/ �/�/�/�/�/�/?"? 4?F?X?C/|?g?�?�? �?�?�?�?�?O0Os/ TOfOxO�O�O�O�O�O �O�O__,_OP_;_ t___�_�_�_�_�_�_ oGO(o:oLo^opo�o �o�o�o�o�o�o�_�_ $H3lW�� ���o�� �2� D�V�h�z��������ΈB�GN_ATC� 1�O� �AT&FV0E�0΋ATDP�/6/9/2/9��ATAΎ,�AT%G1%�B960�+�++3�,.�Hc�,�B�IO_TYPE'  ����Џ�REFPOS1 �1��� x��������?�P� ���6�������V�߯�z���� �9�Ǜ2 1�����$���� �ƿD�ё3 1� ^�p�����:�%�^�ܿS4 1�����Q��Ϻ���q�S5 1��ϚϬ���d�O�|���S6 1�߀/�A�{�������S7 1�����������y��0�S8 1�G�Y�k��#��G����SMASK 1���  
����e�'XNO��;�A������͑MOTE  ���ʔ��_CFG ����<���̒PL_RANG���q���POWER ���^ ��SM_D�RYPRG %��%��dTAR�T �V�
UME_PROs� �ʔ_EXEC_E�NB  =���GSPD� #��4gTDB>PRM_.PMT_m�TQ �����OBOT_N�AME ����׉OB_ORD_NUM ?V���H86�3  �t ���!\<� � # 	r*!�@�"D|<���P�C_TIMEOU�T6 x��S23�2
1�� L�TEACH ?PENDAN_ ����e����M�aintenance Cons�r����*"�/�KC�L/C� :����/? No Usee��/U?�v#�NPO218�����t!CH_Lf� ���7�	�1~�;MAVAIL��a#�������SPA�CE1 2�ٜ �?%dH�9�eF�%�<��L8�?H �9�O�?�O�O _�O(_#WTOfOxO�O 8_�O�O�_�_�__o  i��4mT_f_x_�_ �_�_�_�o�o�ooP .�5;A2@NRO dovo�o6�o�o��@��4��I�N{3] o���S�������ޏ0�Q�8�f�N{4 z�������p��� �8���M�n�U���N{5������͟ߟ��� %�4�U��j���r���N{6��Ưد�����  �B�Q�r�5χϨϏ���N{7ѿ����� ��=�_�nߏ�Rߤ�������N{8�� ��$� 6���Z�|ߋ��o����������N{G �N�� ���$
�� C�e#p����� ��������:hL���2� �+��^�!dt Y� k������� ��8oR~q ������// =/7Ikm�/� ��/�/�/??+?=?�3/]?W/i/�/�= `�� @NP�5< �?�/�) A�5�?1O COI?#J$OVO�O�O�O ~O�O�O_�O�O�O_ ^_ _2_D_v_�_�_�_ �_�_o$o�_�_
o<o�~o@oN<
O�oN{_MODE  +�^�iS �+��ox?v:_��?'y�z�	��o�CWOR�K_AD�mvϽ�q�R  +������p_INT�VAL�`@�zR_OPTION1�� u��VAT_GRP 2�+�w]�(���L��ԏ揥� 
��.�@���d�v��� O�o���dX�ß��� �ϟ1�C�U�g�)��� ������ӯ�{�	�� -���c�u���I��� ��Ͽ��ϛ��;� M�_�!σϕϧϹ�{� ������%�7���[� m��Aߏߵ����ߛ� ���!�3�E�W���{� ����s�������� ��/�A�S�e�w���� ����������+ ��Oas���? ����'9K�[����e�$�SCAN_TIM��a��\��R ��(�30(�L}8z��p%�p
WtZ��2#Nq!�#Y�:.(/1+�#M"2{$!"!d�(~!�!�r #])�0��/�/�/�rܪ)�/  P5:�0�2  8�?xU?g?>1D��j? �?�?�?�?�?�?�?O�#O5OGO?Nq�%ARO�O�O[N![q�;�o�t�Nqp�]M�t��D�i�t!c{  � lM"Nq�A!
%�1_ C_U_g_y_�_�_�_�_ �_�_�_	oo-o?oQo couo�o�o�o�gS�o �o�o'9K] o������� ��#�5�G�Y��o�o �K������Џ��� �*�<�N�`�r����� ����̟ޟ����1�  0�B|�_g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ�p��� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑ��ϐ� ��������0�B�T� f�x���������� ����,�>�P�J�V�  �1���������� ������1CU gy�������	 �y3" HZl~�������C&5/</v+&�r! 5/�q-	12345�678R���L{0�@�/�/�/�/�/?3,?>? P?b?t?�?�?�?�?�? �?'OO(O:OLO^O pO�O�O�O�O�O�?�O  __$_6_H_Z_l_~_ �_�_�_�O�_�_�_o  o2oDoVohozo�o�_ �o�o�o�o�o
. @Rdv�o��� �����*�<�N� `����������̏ޏ ����&�8�g�\�n� ��������ȟڟ����"�+&s�C�U�:��Z��������Cz�  Bp   ����2/$@��$�SCR_GRP �1�(�e@(�l�� �@ Z! �U!m�	 #�-�=�6� n�p�l�S�y(J�w�e�ܞ����3%Dʰ֠o��ป���M-10iAo 890�%90� �Ɓ M61C ��#�-I���#�
\�l�,�O'|�Z!�S�;�o�}�	n�������h����X �,� ��Y"N�a����ߖ�i� @�.!`/��m�����"�.�B�Š�J�H��a�H�A֠p�  @. ��l��?���D��HŠ���H�F@ F�`������ �;�&�K�q�\����� ��<�����������B���YD} h������� 
CҾ?4#��0/v/�%��
��������V�j�@�܆�/ B�*'���P���EL_D�EFAULT  �C�����X!MIPOWERFL  P�xp%W"} WFDOe&� p%��ERVE�NT 1����I�n#=�L!D?UM_EIP��(��j!AF_I�NEd ?�!FIT�/7>�/[?!K�΀? �J?�?!�RPC_MAINĨ?�8��?�?�3VI�S�?�9��??O!�TP2@PU6O�)d�.O�O!
PMON?_PROXY�O�&AezO�ORB�O�-f�O�#_!RDM_S�R��*g_o_!�RL(�_�$h^_�_!%
�0M�O�,i�_o�!RLSYNC�o.i8�_So!gROS�/zl�4Bo �on?�o2S�o�o�o �o5�oY }D� hz�����1� C�
�g�.���R����'�ICE_KL ?�%�+ (%S?VCPRG1��������3$�)��4L�Q��5t�y��6�����7ğɟ�H=��/�9��� �_A���i����� �>����f��끎� 	�끶�1��ޟY�� ����.����W�ѿ �������!��ϯ I����q������ G����o������� ���9�;�翹�˂� ҏ䀄���á������ � �9�$�]�H��� ~�����������#� �5�Y�D�}�h����� ����������
C .gR�v��� ��	�-Qc N�r�������/)//M/��_D�EV �)��MC:U(��]]g$OUTYB`!�x&c(REC 1����` �  ` � 	 ` ` ` ` �!�!U+�#��IU/�.�$1�"T?`!` 8:�
 �P�b6� s�'�  ��  '� �/  =0f���"T�#�!� ` /` ��` ��=y �y �y �����` B�� D�?O�%��|0�ހ<S  ��H�� �0_��? VO�` �4)` M��?��`!y ��0�` k� NPO�OO+c݀;[0�0�1�o  �� iV�O !� � �04�,` �xO��y ��!�Dn� M�O]_�OKc��O�@�F��O�
__._@_R_d_If_�6r _�H�i@U�4�x�C�@��_��!r` �` C` ��P#�_�fy �*y �y �y �<1To�ooh$0k � � � �1   +�i@=�o ;@�2l�0�   K`$|o+�dy �y �y Dqa��! a�oh[�l��0k`�bR  EȢ lP
5�2` ��` �(�c�4�D��!��t~�j��0k� ��3}��`  #"��j2;� ` L` �\� wO���y �y 	��qy ��QX���tkaĀ<Đ?g����?�?�?�?��ď"F V�;T�f�4���R'�+�` =� �� ���
` Q� ,��U����H��` U� F���x�02y0 � � T�B�x�f�������ү ������,��P�>� t���h�����ο��޿ ��(�
�8�^�Lς� pϦϔ����Ͼ� ��� $��4�Z�H�~�`�r� �ߢ��������� �2� �V�D�f�h�z��� ������
���.��R� @�b���j��������� ����*<`N��r�����%V7 1��, P 8� �:���*��o �
Z�!Kd'TYP�E�/e"HELL_�CFG���&� ���"�� %RS �p���//?/*/ c/N/�/r/�/�/�/�/��/?�/)?8;�p:>����` %K?y?�?F=J1J1�p gA�=�1��p��a22!�d��?�?�HK 1���a�?AO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_~|OMM ����_FTOV_E�NO�nwOW_?REG_UI�__?IMWAIT�Rq\�6kOUTf� iTIMe���ZoVAw�1o#a_U�NIT�S�fwMO�N_ALIAS �?e�Y ( heH�o,:z�o ]o��>��� ���#�5�G�Y�k� �������ŏ׏���� ��1�܏B�g�y��� ��H���ӟ���	��� -�?�Q�c�u� ����� ��ϯᯌ���)�;� �_�q�������R�˿ ݿ��Ͼ�7�I�[� m��*ϣϵ����τ� ���!�3�E���i�{� �ߟ߱�\�������� ���A�S�e�w��4� ����������+� =�O���s��������� f�����'��K ]o�,���� ��#5GY }����p�� //1/�U/g/y/�/ 6/�/�/�/�/�/�/? -???Q?c??�?�?�? �?�?z?�?OO)O�? :O_OqO�O�O@O�O�O �O�O_�O%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3o�_Woio{o �o�oJo�o�o�o�o��c�$SMON_�DEFPRO ����4q� *SY�STEM* . �"vRECALL� ?}4y ( ��}6copy �md:progr�am_1.tp �virt:\te�mp\=>des�ktop-b25�t4o0:836?0  916����z} xyzr?ate 61��r@��8�J�\��q
�w ��"���ŏ׏��0:544����6�H�Z��1���!��� ğ֟i�s�����:� L�^����'���ʯ�ܯo�:��frs:�orderfil�.dat�mpback���/�A�S��f�1��b:*.*	��0 &���ɿۿ6n�5x��:\}����������;�M�_�}6��a��Ϝ�,Ͻ��� ������*�;�M�_� r�ߖ�(߹������ �ϐ�&�7�I�[�n��� �ϵ��������χ� "�3�E�W�j�|���� ���������ߍ��/ ASf�x�	��`� ��������=O b�t���*��� ����(9/K/]/p //��/�/�/n�/@�/�/4?F?X?k�!t�~��15432 ? (?�?�?�?p9|��?�?1OCOUOh�7���O2 ,O�O�O�?t?O _�O;_M___�?_�_ (_�_�_�_pO�O~_�_ 7oIo[o�Oo�_$o�o �o�ol_~o�o�o3E W�_�_o ��� �ozo�/�A�S��
;�������ӏ�
2t�����8�J� \�o*}/?�+���Οa�7t/����*���>� P�c�u��������ί a�󏎯���:�L�^�� �$SNPX_�ASG 1�������� P 0 '�%R[1]@1�.1`���?��% ��ֿ����ݿ�0�� :�f�Iϊ�m���ϣ� ����������P�3� Z߆�iߪߍߟ����� �����:��/�p�S� z������� ��� 
�6��Z�=�O���s� ������������  *V9z]o�� ���
��@# JvY�}��� �/�*///`/C/ j/�/y/�/�/�/�/�/ �/&?	?J?-???�?c? �?�?�?�?�?�?O�? OFO)OjOMO_O�O�O �O�O�O�O�O�O0__ :_f_I_�_m__�_�_ �_�_�_o�_oPo3o Zo�oio�o�o�o�o�o �o�o:/pS z����� �� 
�6��Z�=�O���s� ��Ə���͏ߏ �� *�V�9�z�]�o����� ���ɟ
����@�#��J�v�Y�r�PARAoM ����_ �	�z�P���j�OFT_�KB_CFG  �����ѤPIN_�SIM  ��Ʀ�)�;�ɠr�RV�QSTP_DSB� �Ƣw�����SR� ��� & �������ΦTO�P_ON_ERR�  ����P_TN ���AݲRIN�G_PRM� ���VDT_GRP� 1����  	ʧ��\�nπϒϤ� ����������%�"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�w�t� �������������� =:L^p�� ���� $ 6HZl~��� ����/ /2/D/ V/h/�/�/�/�/�/�/ �/�/
??.?U?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o Fomojo|o�o�o�o�o��o�o�o30ѣV�PRG_COUN�T����^rENB)�YuM�s㤐_UPD 1��8  
G��� ��'�"�4�F�o�j� |�������ď֏���� ��G�B�T�f����� ����ןҟ����� ,�>�g�b�t������� ��ί�����?�:� L�^���������Ͽʿ ܿ���$�6�_�Z� l�~ϧϢϴ��������VuYSDEBUG�hp�p���d�y�S�P_PASShu�B?.�LOG ���u�s������  ��q��
MC:\Z�
�[�_MPC`��u���ߒ�q��� �q��S_AV �c���l������SV��TEM_TIMEw 1��{ (�p�Ҫt���s�N|T1?SVGUNS�piu�'�u���ASK_OPTIONhp��u�q�q��BCC�FG ��{I� qB��5�`5� ;zC�l�W�i������� ��������2D/ hS�w���� �
�.R=va������� �/��B/-/f/Q/ �/�/�� �/�/�/ �/�/ ??D?2?T?V? h?�?�?�?�?�?�?
O �?O@O.OdORO�OvO �O�O�O�O�O_�H� _,_J_\_n_�O�_�_ �_�_�_�_�_o�_4o "oXoFo|ojo�o�o�o �o�o�o�oB0 Rxf����� ����>�,�b�_ z�������ΏL���� �(��L�^�p�>��� ������ܟʟ�� � 6�$�Z�H�~�l����� ��دƯ��� ��D� 2�T�V�h�����¿x� ڿ�
��.Ϭ�R�@� bψ�vϬϾ��Ϟ��� ����<�*�L�N�`� �߄ߺߨ�������� �8�&�\�J��n�� ����������"�ؿ :�L�j�|�������� ������0��T Bxf����� ��>,bP r������/ �//(/^/L/�/8� �/�/�/�/�/l/? ? "?H?6?l?~?�?^?�? �?�?�?�?�?OO O VODOzOhO�O�O�O�O �O�O�O_
_@_._d_ R_t_v_�_�_�_�_�/ �_o*o<oNo�_ro`o �o�o�o�o�o�o�o 8&\Jln� ������"�� 2�X�F�|�j�����ď ��ԏ֏���B��_ Z�l�������,�ҟ�������,��J��$�TBCSG_GR�P 2����  �J� 
 ?�  u� ��q�����ϯ��˯���)�;�N�U��\�_d, �j�?J��	 HC��8�>�����9�CL � B�m�����z���β\)��Y�  A���B��;��Bl�=�,�����Z�,��  D	 �{�F�`�j�Cs���H�Ϧϰ̖���@J� �+�>�Q��.�|ߙ�@d�v��������؈J��	V3.00~m�	m61c��	*,�$�I�;�D�>���J�(��� qr�D�s�  #�����D���N�J�CFG ��ef� i������������� �7�E��E�k�V��� z��������������� 1U@yd�� �����? *cN`���� ��m����/"/� U/@/e/�/v/�/�/�/ �/�/	??-?�/Q?<? u?`?�?�?J�6��?� �?�?�?*OONO<OrO `O�O�O�O�O�O�O�O __8_&_H_J_\_�_ �_�_�_�_�_�_�_o 4o"oXoFo|o�o���o �obo�o�o�oB 0fTv���~ �����>�P�b� t�.���������̏Ώ ����:�(�^�L��� p�������ܟʟ �� $��4�6�H�~�l��� ��Ư���د�� ��o 8�J�\����z����� ���Կ
���.�@�R� d�"ψ�vϬϚϼ��� ������<�*�`�N� ��rߨߖ߸ߺ���� ��&��J�8�n�\�~� �������������  �"�4�j�X���|��� ��n���������0 TBxf���� ���,P> t���d��� �/(//L/:/p/^/ �/�/�/�/�/�/�/?  ?6?$?Z?H?j?�?~? �?�?�?�?�?�?OO  OVO��nO�O�O<O�O �O�O�O�O_
_@_._ d_v_�_�_X_�_�_�_ �_�_o*o<o�_oro `o�o�o�o�o�o�o�o 8&\J�n �������"� �F�4�V�|�j����� ď������O�$��O ��f�T���x������� �ҟ��,����b� P���t�����ί௚� ����(�^�L��� p�����ʿ��ڿ �� $��H�6�l�Z�|�~� ���ϴ��������2�  �B�h�Vߌ��8��� ��rߠ�����.��R� @�v�d������� �������N�`�r� ��>�������������  J8n\� ������� 4"XFhj|� �����/0/�� H/Z/l//�/�/�/�/ �/�/�/??>?P?b? t?2?�?�?�?�?�?�>�  @
C �
FO
B�$TBJ�OP_GRP 2���5�  ?�
G6B=C��DL��0�xJ�@��
D@ �<� ��@�
D �@@UB	 �C��� �Fb  C�xVGUAUA>����E��E�I>��@�A�33=�CL�@�fff?�@?�ffB�@Q�E-_8W�N���O>�nR�\)�O�@�U����;��hCY�@��  @�@UAB� � A�$_�_�S�UC�  D�A�LwP��RO�z_�Sb���
:���Bl�P��P�D�Q�_So
A?Aə�A�hcZQsDXg�F�=q�e�
o�@�p��b�Q�;�AȰ@�ٙ�@L�CD	�x`�`�o�ojo|o>BÏ\u�oh�Qts}�a@33@QV@C��@�`ew�o>��D�u*�@�� p�qP<{�Nr�@@�PZv_p�� ��&�:�$�2�`��� l�&���ʏ����!� ����@�Z�D�R������DT�
Fґ�E	�V3.00�Cm761c�D*���D�A
�� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,I&�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^'`;Q���8�E`F�O���
F���Q��K�2DES�TPARS  ��8O@3CHRe�AB_LE 1�DK.�
CP�%� ~ �P��P�P�	GAP�	�P�
P�P���
A�P�P�P�|�RDI��NA����¿Կ���`�Oh�z˄� �ϨϺ��΀�Sf�LC *ʍߟ߱������� ����/�A�S�e�w� ���������)Me� iߘ�$���1�C�￀��%�7�IȀ�
�N�UM  �5*NA�@@ ��[����_CFG ������A@6@IMEBF_TTk���LCx�5VERY�6�K�5R 1�DK
' 8�
B@� �0/�  ��� ���� 2D Vhz����� /�
/S/./@/V/d/�v/u_��b@L
�6@MI_CHAN�A L �#DBGLVPCL5A� �ETHERAD �?�550�M���/�/N?0F� ROUmT_ !DJ!�4��?q<SNMASK�*8LC;1255.��5��?�?2DOOL�OFS_DIk���%9ORQCTRL �mK���hM8WO�O�O�O�O�O�O �O
__._@_�|ON_�`_�_a�PE_DE�TAI8-JPON?_SVOFF#O�S�P_MON ��J�2�YSTRT�CHK �DN�g?�RVTCOMP�AT�X53�T�PFP�ROG %DJ%}	qaRAM_17o<�\APLAYl��Z_INST_M�0e �l�W�dUS_�WoibLCK�l�kQ?UICKME� #�ibSCRE@p>-:tps�ib �a[p`y�"qp_uy���Ti9SR_GRP� 1�DI ؕ�0��z�� �5�#�Y�G��2 �� ��S��o����܏ǅ�� ��)��M�;�q�_� ������˟���ݟ���7�%�G�m�	1?234567堃����b�XZu1��{
� �}ipnl�/ՠgen.htm�����*�<�R��Panel _setup@�}6o���������ȿڿ  o�e��$�6�H�Z�l� 㿐�ϴ��������� ߅ϗ�D�V�h�zߌ� ���C�9�����
�� .�@��d��߈��� ������Y�k��*�<� N�`�r��������� ������8��\�n����-�nU�ALRM�`G ?=DK
  � 	L?pc�� �����//6/~�SEV  ��h&�ECFGG ��]�&��A�!�   Bȣd
 7/�c-5�/�/�/? ?%?7?I?[?m??�74t!�r��[ �3ȏ��?B'Imf?wk�P(%*/O`
OCO.OgO RO�OvO�O�O�O�O�O`	_�O-_�<�d �=��?;_I_?pHIS�T 1��Y  �(�  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupage,153,�o��_�_oo �� �_�]936�_lo~o �o�o1b�o�o�o�o %�oI[m� �2�����!� �E�W�i�{������� @�Տ�����/����S�e�w���������� L��QL������1� C�F�g�y��������� P����	��-�?�ί �u���������Ͽ^� ���)�;�M�ܿq� �ϕϧϹ���Z�l�� �%�7�I�[���ߑ� �ߵ�����ğ֟�!� 3�E�W�i�lߍ��� ������v���/�A� S�e�w���������� ������+=Oa s������ �'9K]o� �������� ��5/G/Y/k/}/�/� �/�/�/�/�/?�/1? C?U?g?y?�?�?,?�? �?�?�?	OO�??OQO cOuO�O�O(O�O�O�O �O__)_�OM___q_ �_�_�_6_�_�_�_o o%o/"/[omoo�o �o�o�_�o�o�o! 3�o�oi{��� �R����/�A� �e�w���������N� `�����+�=�O�ޏ s���������͟\�����'�9�K�6o���$UI_PANE�DATA 1�������?  	�}]���`��ȯگ��� ) � $�ᔒ�O�a�s����� ���Ϳ�����'� �K�2�oρ�hϥό������������ Ha$�7�<�N�`�r� �ߖ��Ϻ�-������ �&�8�J��n�U�� y����������"� 	�F�-�j�|�c�������������� +=��a�߅�� ���F�9  ]oV�z�� ���/�5/G/�� ��}/�/�/�/�/�/*/ �/n?1?C?U?g?y? �?�/�?�?�?�?�?	O �?-OOQOcOJO�OnO �O�O�O�OT/f/_)_ ;_M___q_�O�_�_? �_�_�_oo%o�_Io 0omoofo�o�o�o�o �o�o�o!3W> {�O _�_���� ��pA��_e�w��� ������&����܏�  �=�O�6�s�Z���~� ��͟���؟�'�� �]�o���������
� ۯN����#�5�G�Y� k�ү��v�����׿� п���1�C�*�g�N� �ϝτ���4�F���	� �-�?�Qߤ�u߇��� �߽��������l�)� �M�_�F��j��� ����������7��[�����}�l�������������)��$�� Pbt��� �����(L 3p�i������ /(�����$U�I_PANELI�NK 1����  � � ��}1234567890Y/ k/}/�/�/�/�$��W/ �/�/??+?=?�/a?�s?�?�?�?�?S9S h*�=��U   �? O(O:OLO^O�?\1O �O�O�O�O�O�O�O_ (_:_L_^_p__~_�_ �_�_�_�_�_�_$o6o HoZolo~oo�o�o�o �o�o�o�o
2DV hz$�����
�E0,/A�M� /�p�S�������ʏ܏ �� ��$�6��Z�l� O����<�?�����T! ���1�C�U�g�Z3 ��������ǯٯ�z� �!�3�E�W�i��<�� ������C��ÿտ� ���Ϥs5�G�Y�k� }Ϗϡ�0��������� �߮�C�U�g�yߋ� ��,���������	�� -��Q�c�u���� :���������)��� M�_�q���������(� ����~���7I, mb����� ��3ƞ����՟ w��������/ ��,/>/P/b/t/�// �/�/�/�/�/??�� ����^?p?�?�?�?�? ?��?�? OO$O6OHO �?lO~O�O�O�O�OUO �O�O_ _2_D_�Oh_ z_�_�_�_�_�_c_�_ 
oo.o@oRo�_vo�o �o�o�o�o_o�o *<N`���� �������8� J�-�n���c�����ȏ ڏI��m"��F�X� j�|��������/֟� ����0���T�f�x� ������?/?A?�o� �,�>�P�b��o���� ����ο�o���(� :�L�^�p����Ϧϸ� ������}��$�6�H� Z�l��ϐߢߴ����� ���ߋ� �2�D�V�h� z�	����������� g�.���R�d�G��� k������������� ��<N1r�� ��;��&8 J=�n����� �i�/"/4/F/X/ ǯٯ믠/�/�/�/�/ �/?�/0?B?T?f?x? �??�?�?�?�?�?O �?,O>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_#_�_ �_�_�_ oo$o�_Ho Zolo~o�o�o��o�o g�o�o 2Vh K�o���������o�/�/�u���$UI_POST�YPE  �%?� 	e������QUICKMEN  ��d������RESTORE �1ݏ%  ���,�>�b�m]��������� Οq����(�:�ݟ ^�p�������Q���ů ׯI��$�6�H�Z��� ~�������ƿؿ{��� � �2�D��Q�c�u� 翰��������ϛ�� .�@�R�d�߈ߚ߬� ����{υ����s�%� N�`�r���9���� �������&�8�J�\� n��{���������� ��"��FXj| ��C����ނ�SCREր?�ۍu1sc�'�u2G3G4�G5G6G7G8<G��USER).2@T(IksQ�U4�5�6�7��8���NDO_C�FG ޖ�  �&� ��PDAT�E ���None V��S�EUFRAME � ��&!RTOL_ABRT1/���H#ENBR/C(G�RP 1���?Cz  A��#�!���/�/�/�/�/ 6
??A*ՀUr(A!a+?MSK  u%}1�a+N.!%[�~2%���?��VISCA�ND_MAXs5�I�](�0FAILO_IMGs0`����#}(�0IMREG�NUMs7
�;BS�IZs3&����,CONTMOU4Q u4��PE�_�c�� �@��"�FR:\�? �� MC:�\RC\LOG�FB@� !�?�O�A��O_�z �MCV�O�CUDM1*VEX3[�`�TqF�"ᖉ�`(��o=��͍_��Z �_�_�_�_�_�_�_o o,o>oPoboto�o�;_PO64_9C�B Κ�n6�eK LI�A�j�h�aV��l�f@�g�o� =	��hSZV�n�����gWAI�o�4ST�AT �+�@�O���z$���5�J!2DWP  ��P G)����a��;@'��2_JMP�ERR 1㖋
�  ��2345678901|����� ��ď��ɏ���� B�5�f�Y�k����<N0MLOW{~�@�0�@g_TIYH�'�0�MPHASE  �%���3SH�IFTO21"x[
 <���?\��;� a���q���Я����� ݯ��N�%�7���[� m�������ɿ�ٿ뿀8��!�n�E������*	VSFT1֝cV�0M�� ��5�q� � ��EA_�  B8����E�� p�����ª�ÌB ��ME$�u4�����a{~&%��M���x[�p�30�$�xpTDINEND]H^8t�Or0U?��[J¨�S�ߏ���s5����Gy�	��,��������ߍ�REL�E �s/q�XOjFt�_ACTIV��~8��
 A �;}�<����RD�`��C!Y?BOX ����V�v��p2��>��190.0.���83����254�����`��� �q�r�obot�ę�   pHa�upc���u���p��r���ZA+BC�#�-,u�  �r�5X?Qc u�����/� 0//)/f/�Z;D�q���