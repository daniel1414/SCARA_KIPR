��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
FPCOU�PLED1 $�[PP_PROC�ES0 � �1z��UREQ1� � $SO{FT; T_ID��TOTAL_EQf� $,NO/�PS_SPI_I�NDE��$DX��SCREEN_�NAME ^�SIGNj�|�&PK_FI� �	$THKYޠPANE7 � 	$DUMMY�12� �3�4���ARG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 � ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4C_WA�4�12HG�W~0�$	Y $D�B� � COMqWƻMOJWH.
� \�VE�1$qF �A�$O���D�B�CTMP1_5F�E2�G1_�3�B��2(GX_D�#� d $CA�RD_EXIST��$FSSB_�TYPitAHKBgD_S�B�1AGN �G� $SL?OT_NUMZIQ�PREV��� ��1_EDIT�1 � h1G�=H0S?@f%$�EPY$OP�c �0LETE�_OKRUS�P7_CRQ$�4�V�AZ0LACIw�Y1�R@Pk �1w@ME=NP$D�V�Q��P��A��G BLv*OUyR ,lA��0V1AB0~ O�L]eR"2CAM_�;1 x�f$ATTR�MP0�ANN�@�IMG?_HEIGHQ�c�WIDTH�VT�C�U�0F_ASwPECQ$M@gEXP;�@AX�f��CFT X O$GR� � S!1z�@B`NFLI�`<t
UIREs3��tGITCH~C�`N�.0S�d_L�`�CL�"�`EDkp;tL0J*DS�0>0�zra�!�hp;G0 � 
$WARNM'@�f�+P� �s�pNS=T� CORN��1�FLTR�uTRA�T@0T�p  $ACC�1
� ���ORI	`!S<{�RTq0_S�Bs��CHGI1� [ Tpu3I�8�TYVD+P*2 ��`v@� 1R*HED�cJ* ���2��U3��4��5��6��U7��8��9��qO�$ <� #p5x�s1v`O_M�@��C t 0E�v�NG��ABA � �c��YQ������@B������P�0X����x�p�P@yP�2� ����J�S_R��BC�J�L�2�JVP�CR�`�}@w��u�tP_}0sOF� 2  @� �RO_����aIT<8C��NOM_�0�1�åq3���T !�#���@xP��J}CEX�G�0� .�<�p�
$TF`��Co$MD3��TO�3�&@U=0�� R�H�2�C1{�E͡� vE�uF�uF�F�0CPo@�a� 	P$@`PU�3�f�)"��)�AXd 1rDU6�$AI�3�BUFVnPȲ�!c |�pڶ�pPI���PZ�MY�M�f�̰i�FZ�SIMQS��/��A-���9��kw Tp{z�M��P�B�FAC5TqbGPEW6���Ҡ��v��MCc�5 �$}1JB�p;�}1DECGڙ�G�F�-�b� ě0CH�NS_EMP��#$GO���+P_��q3d�p�@Pۤ��TC�� {r��q0�s��a�/�� `�B���!	���JR!0���SEGFR��ITv �aR�TjpN%S.+�PVF�����ʹY�K��a1��)B���( ' j�Av�u�ct��aD�.0����*�LQ��D�SI!ZC������T��O������aRSINF �����jq��C��C�����LW�����x�C3RCLuFCCCkpy� ����N}���bA��������d��DwIC��C���r��+ P��Lz�2EV2�zFH�_��FpNt/��>����H�1Q��!  ��@�Qx ����U�kp�2 ��a��s�+���qRT!x "�4�4u2���tAR���`CW�$LG�p��B�1�Pr�P�t�aA?@z�ϣ~01R�ӲME�`8�oC�RAs3�A�Z����pb�OS�FC�b�`�`FMp�� �0��ADIS+�aV% ��b�z��pE$�pRp��cV�S�P��a+QMIP5�`Y8C��MeҰpU��aUS" ]$=�TIT�1�S��SG1��#�8��DBOPXWO! T#���$SK��2��D�BTmTRLS$�l�Q0TQ��P`P�D��q�1LAY_CA�L�1�R^0o f7PL)A�Q�D'a�73a�7���o�DB!S%�2?�PRj� 
p*0���S& =�6A$��$ �*ЅL�9'�?'�U�T(�ODCS)#ODE3NE��*BO'��0RE�pB+H� �Ou�&$L�C'$�3R��K42�LVO�_D~!U�ROSbrq�v�R���~�CRIGGER�F�PA�S��6�ETUsRN�B�cMR_}��TUbp���@EW5M$���GN=`����BLA��TUܡ({$P�)$P "s�*hP3a��C�TΣ@DO>���D�A����FGO_AWAYF�BMO"�a�!*0wCS_P,<aISt�� �� �s�S#�Q���Rw�c�V��Qw2�VW��'dNTV(��RV;���� ~��mgŃ��Jt��<<@��SAFEڥ�f�_SV�bEXCL�UT��� ONLď��cYfЀ�y�OT=EuHI_V} ��PPLY_�q7�VRFY_b3���Rj L�_ -h@0��9_y�1� J�Q;SG�  .�rŐ 1PNQ5�� _q���;P☐Vby|rsvANNcUN<@�$�tIDX�	UR�c[P� �y�q�i �z�vIrEF�PI:<B/��$F�r�$�АOTQP�A ?$DUMMY��&����&���*0t�U0o `  �HE��\���^r�cYRr SU7FFI���Pa0(��P)�5#�6#���DMSW�U1 8� �KEYI��4�T�M�A��ځ3QՆIN�ݱv�4:�Dj P2{ D��HOST�0!�������������EM&����n*0SBL� UL��3 Z���D�)1�T�@S4 � y$���USAMPa�@��.������V I�@|��$SUB�����;@c����3��SAV���������X��`�vP$�@EC!�	0YN_B35 M0�pDI�t�PO\��M��#$E�R_I�B� �ENC2_S�T6X��2������ �cG���0 BS72��1��A��>��8  ������@PK�Dk!uq��AVERҁ�����gDSP�ܢPC?����26�\�����VA�LU�HE �M�_�IP(�ܣOPP� 5�TH��ͫ"��S` 4�.�FB�6ad��~�� 5�SC?q����ET�9�ȂFULL_DU ���qKP�ԝ������OT�"T�PNOA�UTOS:�$�YĪ�Z� ���X�Cʮ0h�CE26
�p�V�L� ;H *h�L� ������$P��wc�ě1 �Ʃ1��C��Ƨ��Ʋ����7��8��9��0T����1��1��1	�U1�1#�10�1=ڕ1J�2X�2����2���2	�2�2#�2�0�2=�2J�3X�3R��3����3	�3�U3#�30�3=�3J�e4X�#���SE�2< <8�Z�����I��e�$�}�"qFE85P?PT= ,f��a�? �P�?(i��e�i�E�Pq�Ю1aT>F�$�TP$!$VARqI����UP21p3? 7���TD��s���p��������_B;AC2@ T�����$uP�*��Þ0� IFIw�0�P� � )PB"JF0P�TAt ;u�"�"pu STvt: �b�t�@�l�6	sC2	>0���S����/bF��FORC�EUPsr��FLUS�pHfNn���^�bD_CM�PEv*IN_t�e`.�REM� F�a�@a�0�Te�Kd9N~�eEFF�j�PINJa�OVM�OVA�TRO�V��DT	��DTMX,A��P*���0M(xR#�0�CL*_��u*�Pr�{_XЉ_T�+Xѕ�PASaD% ���(װ�1`�&_A@R�Q�LIMIT_��4�� M��CL�tˑRIVW�*2�EAR�IOxP�C�P���B�R�C�MQP*�b !GgCLF�#�1DY�8�} �q�35T�%DG����0�5N�SSt0��B P��1�A���`_�1�8�11R��E�C�13 K5 FO�GRA��gC��ik�`W�ON��"EBUGwctBx�#pC ��_E D� �� q �T�ERM�EE�F#pO�RIS�@F�Eא�GSM_�`���@G�E�q��TA�IH�IU}P��I� -�QƯ�D|`�C|PE$gSEG#Z�0EL�ewUSE�PNFIz�LRT�kA,��DTF�$UF�`O�$\��a�P/���Wi@qT��t �cNSTT�PAT��h��RPTHJKa-�E
�65MR�<p&�WUw�&�Q�LQRx<`�Y�qSHFT���MQ�Q�X_SHOR(�*��F �@$�GM`9H�u OVRq��qR6`I`4U� �a�AYLO���"J�I�u2b��Q��oƸ�ERV���a� 6j�WnP@�R~�E �e��E Rb1=Pp�ASYM|�p�FMQWJ`W�� E���Qy�b0�U7tnPI��Uw�/�ePo��`o��fgORnPM��G@SMTfJg�G1R��aC�qPA|P���p=��K � :FTOCFQ�yP9`N $OP@�/��#��N �!O,�ڐRE
�RdS�Q�O����Re�R�UN�%�a#e$P�WR0IM@��bR�_ ���=�mR L�VBH�_ADD�R$�H_LENG��Rǁ���T�R� S.O�M H�S��恀~�������	�S�E!u���S:�MN�1N��p��F¹�OL��8�3�x3�=��ACROc� z�P$��[·a;� N �OUP���r_�I���q�q1�ѭʓ ��ԙX!՘Y1՘t!՘`	�ԙлE"IO����DϗA�ߕ9�g�O $���p)_O�FFb�;�PRM_�Ò_HTTP_�[�HjP (��OcBJ�2��#$$��LE�S���Q � ���AB_�!T���S�p;x �LV��KR32@�H�ITCOUBGE�LOہ磴!��`@��"�G#�SS�F�HWD�SQjR�}lpINCPU4BVISIO���������
������	� ��IOLNS�z 0C$SL�r�@PUT_�	$@��PV0�ɱ)�F_AS�2T �$L  �� =a0U�@9`dQٵ��䳊`�HY#�]�6�_�U9O�3U `"�{��$�5"M�5 Tƥ�R�P�;@��ǿ�T��µ�1�	PJeV]���N�EfgJOG{W��DIS��K��� �3W XХQVv��P;��CTR�S:�FLA�GBB�LG�tX ��� ���aCLG_SIZ����d ��,���FD��I�ا� ��׏ث@�֎���� 	�d 	��	��	�@<	�% SCH_��R�H��aBg�Nє�Y��!E�2��p�J �U}�}��pL��|�DAU��EA�����t����GH�r_%�B�OOZh A<�f0IT2���@8�wREC�SCRB��=�D:�����MARG�<18��0��Ha�%�Sȣ$�W?��%���0�JGM��M�NCHz%�FNK�EY��K��PRGƾ�UF��g`��FW�D��HL	STP���V��mP������RES;	Hp��-�Cid@6r0�.0s��	U|����r�Xb��P�E���G��`PO�
.��M�FOCU�RwGEX,�TUI��	I��p�K|�V�� V����A`B���p��A`�Nu��SANAx%�FR��VAILy��CLP1uDCS_CHIyD�
��O�DX1�S� ��S�V�IGN��~�ӽ��\�T���_BUFUF�1[5�o`T�$��� ����B���*A��\5�o`ܰ���c��pOS1�%2��%3�!�A��0] � ܩ�qEU��\���IDX�tP�b�D�O� ��Q6ST�|�R��YV�@1 /\$EO6CO;��{�^6q6�&��0^ L��K�[@`�9`(���S���:�����x��_ _ o�p�ÐЌ�� C�@Cp�` =�� CLDP|�uTRQLI��Ft
�4I"DFLGV�"@1�VC�D)�VGr�LD8VE@DVEORG
�q iB_�g�H
��d�D�ta �M�@Dr1D
VES�pT4@I��@T}VRCLMC%T`�O�O7Y��0MI�έtb dy��!RQzI�M�DSTB��0 �VO�XAX�r �X�\EXC+ES6�sUM_��qc6��Rt��vR<�j�pd��V_A�Z���(k�_�X@K�te� \����/�$MB�s�LI���cREQUIR�b��l���h�DEBU����ML
�0M,�f�r=��`��4��%RsQND���p±pgw�n�?�sDC��IN����p�,x' NV���K��R� qPST� hn��LOC�&RI���%EX�vÀ�!�Q�sQODAQ,�i �X��ON���MF \����v9�2%��5�u�k�0���FX�PIG}G�� j �M�@�2!���3��4R �%?3;�|�K�|�Z�<G`E�DATA{'��AE�U��1!በNZ"�k t $MD
��I��)Ɔ ф��фH�p�`Ѕ�X�҃ANSWe�ф�!'
хD[�)�r��P���l �PCU��V��X@�uRR2��m� D���a���Rd$OCALI�P"�G�:w�2��RIN��z��<u�NTEڰ�"n�I���°r��ڰ_N��oÕޒi�oT۔b�p�DIVmVDH��Pݐ��q� $V؄�+s1$��$AZ�"��� �"f�_��e�rH �$B�ELT>��1ACC�EL!������ICRC��P��t�T31�h�$PS�P'BL�0M�ʤ<C������<���PATH���D���3ТZ��Q_�! U�2�8�R� C堌��_MGP�$DDxU���/�$FWh������q�����f�DE���PPABNاR?OTSPEEH��!��4@J��!��P��~�0$USE_��2�P��O�SY��g�ZQ B�YNyPAO���OFF��MO�UR�NG�O�OL�L�INC.��q���u��Rn�PP�RENCS�����Rȡ���TŠIN'2IТ���`R��VES�{���23�_UPI���LOWL!� �4@���D� �R{`���0��5b9Cΐ��MOS4 Ld�MO���PWPERoCH   �OV� �b��!m�@1�^T@1��s��hP�`�� V5�'`ѡ��L���Ig����UP�Ӛ����TRKv�#2AYLOAA��$a1�Т@�p5�p40��RTI(a|�40MO����R$b �@N��T��w�L����"f�DUM2,�S�_BCKLSH_CТ��B�A�u�'�Y�������6�x�aQCLALz ���Ar�`��CHK4@+5SH�RTYS��}%�A��9_:36�_UM(`n�9C{�c�SCL��ʰ�LMT_J1_LDS��P������E������������SP�C��;���	��PC�sѦ�H�0�`Y�q�C�3P�2XTc�g�CNE_��N��i��SH ���V	�*3�Ň�=�Т�AC� y�SH :3��g��ƝA���s�`4�ѡ��c�PAx�&l�_Pw�[�_5@���8�V�4AH�ZK�JG�G"M��OG[��ToORQU��ON.ـQ靰wbLҠᝰ�_	W��1�_A��G��TM��I�I�IM�	F�p�JPQ2(�A_��VC��0�T�RS"1�Y.�Pm/�R`%JRK�Y,�"�&PDBL_�SMh�RM)p_D9LG�RGRV��$0G��$M��!H_ �#�:COS;`�8LN� ;;\%B4G�=9�M�=9!y:g<-!�%Z60L־!MYD1�8$2�TH*=�9THET=0�NK23M�BlA�E0CBFCBA�C�Q�R,B$:AG�:A�FSBG�XBEGT	SaʱC��qW4�&�Dg3�Gv3$DUH�Ih�Aw�x��R�F���QQ���v$NEd�IF0Y�`R�E��	$%��1A�5#U,W
581LPH(eR��RS\%tSg5tSv5R��6�S�Z�6%�VEXV�:X7�]\VlZVy[V��[V�[V�[V�[V�YHEX^Vdb\]�{h�y[H�[H�[H�[H��[H�YO6\OEXOT�i[^OlZOy[O�[UO�[O�[O�[O�6�FR'A�yg5�t8WS�PBALANCE�_�1�sLEo@H_�5SP��X6�rg6�r>v6PFULC�x���w�v5Ț1n}�U�TO_C�nT1T2G���2N*�z��� g���k���@ע�����T��O����IN�SEGz�%�REV8��%���DIF�홳1o҇�1p�@OaBȁ��#��MI���5��$LCHWAṞ���AB*y�$MECH0A�0>�D�Y�AX>�P��]�W(�<�q 
^����n��ROBV�CR��정R1d�SK_|�pj�s P R�_��R��H�Ҕ��1���ԲҐ����Ґ�&�IN���MT�COM_CD n�t�  P�ڀ���$NORE��9����(�u 8�G�R�I�SD�@AB�J�$XYZ_D�A9Q���DEBU���M��U�v �p$��COD�� 褢o�J�j�$B�UFINDX԰ܻ���MORœw $1�U��-��v�LF��� Ң�Gܢ�x � $SIMULX�����$����OBJE�p$�A�DJUSB�5�AY_Io��Dc����nG�_FIJ�=�T����������������Հ�P��D�F�RI��׵T��RO����E����O�PWO� ɐy0>��SYSBU�PΠ$SOP���#�'�yU&�ՀPRUN�M�PA�DL�H�!�.��_OU�!A����r�$��IMAG���ϐ�@P��IM�����IN� u£�RGOVRḎ>°��P����԰�@L_`:����m� RB� ��@M��EDTՠJ� ��NpM.����ETI���SL��pɐz x $�OVSL��SDI��DEXqk�i�=!H{��Ѕ�V���N�р�{��Њӟךط�M��!uG�_SsET�ɐ{ @����g���RI&���
��_4A��	����ׁ|@��  | Hϑ�I�J�ATUS��$TRC�@ǰˢD�BTMM�7�Ij����4��#�,�ɐ} �DϐE~�k�A�`E�ۂBᏱ
��B�EXEH�Z�ќ��{���1~��АG�UP���s$����XNNm��=!p�L!p� �PGn&��!UB6��g��6�
�JMPW�AI� P��N�LO��j�F��#�$R�CVFAIL_C�j�Q�R��Q�Z�M�� 𣕠���0R_P=L
�DBTBm��j�BWD��A�UM���IGe���m�� GTNL� ����R�D��.�Ep����DEFSPy� G� Lϐd�7 _: H�HUNI��r�F b��R��^�� _L��5P@����P�ȑ����F����Ѐ��p:��N�pKET�}��� P��ȑ� h~W�ARSIZE���l���S@�OR~
�FORMAT3����COJ����EM2V�lUX�����PLI��ȑ� � $#�P_S�WI��բ ����A�L_ ��E AR��B�,@C��Dj��$E���uC�_��	� � �c ���qJ3�@�����TIA4�5:�6��MOM��������#�Be�A�D�&�&�PU;@NR�J%�J%��EŔ�� A$PI�F�ޑ��$ �%�#�%�#�%=D�&�+ QD�DpсF���U�|��g�SPEED�`Gd*4f�7167f� ��16g3@8��O9��f�SAM�p맣417�3f�MOV���D�1@ƀ�E�4�E�17 1��42�������5n2��Hm��3IN2Ln �39HUK0Df�;J{HRD<{K�KGAMM�v�A>�$GET��Ƞ�L�D� �
b�LI�BR��I��$H�I��_��P��bVEĂXA^:P+VLW ]XVO\:Y|V+V�V������ $�PDCK�U�L�_�0�� �.B�m!E��W��T&�Yr ��$I�RS�D`��&����(�LE�`ޑ�Oh�)`� ���H�ɐ�P��UR_SCR��a^���S_SAVE_�D�īe��NO�C ����`�D��&�i ��)�iapz{p�� �&Ex@�q��0�B�� �5G�2�+8!�;6�� g8�w�ucs�1����HM{%� ����!G ����c�w���`ζ�q!W�`��$��0�N ���R�qM��H�CL�G�GM�aǒ� �� $PYr�3$Ww�+�NGt�� w��u��u��u���������@[L�nX� O�mZ��GQ��Ŕ� pW�#�c �&�o�o#5��_)�� |Wи�` ��������`�ޗɖ�EQ��EB���b��� ���P���PM��QU�0 �� 8� QCOU�as�QTH��HO�L��QHYSES�1[�UEG��b� ]OM�  �P4��U�UNI�J� ��O��)�� P��������a��ROQG�j��2��O��c�󠉠INFO(�� ��ث�
��ȏOI�� (`SLEQ"6D�5�D�ܦ����DS𿠒D��VPO�P�0#3Q�EMPNU����AUyT�a��COPY�1P�಼��`M��N�������CT�� �R�GADJ(���X#�_$� '��'�W%�P%�]`'�:3��;�EX��YC��$�@OՐ(���7_NA�1!S����i����M� �s ��p�POR��Ì&��SRV��)l����DIT_p� �� ��
��
�w�
�U5�6�7�8��ҏS�b�����MCS_Fe��pL�a�a{;�Rq���/���җ#�0��k��� �,`FL����`Y�N{���Mp�C��GPWR��������ODELA �6Y��ADR��QSK;IP{%� �����-OŀNT�1�0*�P_����I�`߂̐ `��#`�3`��n�k n�;�m�H�m�U�m�b�zm�98a�J2R.0n��� 4� EX�@TQ����q����������y`RDCNx�� ���X��RF�E@AY�_�X�D�RGEAR_�@I9O�t=bFLG����EPC��UM�_���J2TH2yN�# � 1�U�A�G�@T�P �$"���M��-�I���4��REF�11(��� l!�ENAB� ��TPE2`{�  8Wܠ�M�q�CL@��R�w��2'�-?Qcu��3'�������4'�'9K�]o�$�5'���������6'�!/3/E/W/i/{/
�7'��/�/�/�/(�/�/�8'�?-?�??Q?c?u?�SMS�K(����� E��a�REMOTE���
��`/B`�L�q-CIO�UQEI�0��R� W\`��� /���-�%� �ӿ����ՈB$DSB_SIGN'a�q�����C��pS23�23E���$�DEVICEUSKC�r�r�PARIT!�AO�PBIT�q��O?WCONTR���qX�0�rCUPM�s�UXTASK�SNxq��P�DTATU�p!�P�A3`���u�e��_�pC��$FREEFROMS�������GETA`��U�PD��AEbSP|TP���� !�8$USA�����9<h�{�ERIO���`&ՐRY�U�B_�`��qP�QQfWRK�?��<Dh�3fh��6FR�IEND�qg�$�UF�U�p`TOO�LwfMYd�$L�ENGTH_VT�ߤFIR��cM�SyE�@�iUFINtr:аARGIaF�OAITIi�gXF�l�i�fG2�WG1��0 �Sr$wPR��sa�u�O_�@�P��xQR�E���SU�ءTCp�N�=qyv �G��]R���u��Q�A�� hzhZUz�ZU�t���|{P�T�X �P*��L��TcH��hPh�U�T�SG��WX�)��r>�D���.���C�z�N�b��$�v 2�!�-a' R3i1?h.`21k2��31k3?j���@i�����6{��s{��r$V��bV�eV���vYr
���O�[V{�@���hv3Ru�^pib��PS��E�$���c��5$A8й�PR)��u,�S���@��� �A�R�¯ 0�p�v���P�N�����!��P>p ��
�US^zA� �\�R���GA_�Š��Ny@A)XQ��Ag`L�ag�^p�THIC'a��8-����QTFE���>m�IF_CH'cp�aI_����6D�G1՘�٤*��h��`��_�JF�PRW�I���RVATF�� ��\�'�f`��)�DO��e)�COUW�C�A�XI�D�OFFS=EZ�TRIG�sz��,�)�#g���z�Hx����g�IGMA�P��a\���ȸORG�_UNEV#@Ͳ ��SD���d ӎ$����GR3OU[A�TOa�Q��DSP#�JOG�V�S8�_PV�3RO����U�mpEVKEPF��IR?�_�=pM �&��AP���E�������SYSv��B��;PG��BRKYr����b�\���������k�ADVQ�y�BS�OC�C@N�DU�MMY14��`S}V�DE_OP1S�SFSPD_OVR���C~�N�QÓOR\׶0N�P]�Fء�]�<�OV?�SF��a����F���Ac��As�؁a�BLCHD}L�RECOVM��P<�W�`M<��?�#RO1S�K�_a�_�� @���`VER�t�$OFS�`CV�@_bWDv� �rѰ��R��9�TR%Q|A�E_FDO�ƟMB_CM[A��B/�BLl�_¦�l�甁V�qDb�P����G���AM�Ú�yP��'��_M��>R��HC4�8$CA2���Ȱ>��8$HBK�Q��N�IO1e]�iAA�PPAQ�}�b���u���iB4�DVC_DB�c�񓡦B����A"��1��'���3��-�/ATIO�@��FP�M�UDc1�HFCAB H�0bFs�p�p��Ea�<�_BP��SUBCPUk�I�S%��@�� ��P�s�,���B��?$HW_C!���i��x�A'q\�l$�UNIT��l�A�T}����I�CYC=L��NECA#���FLTR_2_F�IҤ�H)�FEaLPxU˲���_SCTosF_�F��
v�
�FS�A���CHA�Ja^���3R�RS�D1�B ё�l�i@_T��PRO ~�)PKEM�0_���8��3� �<�*%D�I�P��RAILAiC��rM��LO��c+�i���-��-V'�PR��S{q*�ҕ!C���@	&�FUsNC�³�RIN�p`Z�+`? �$(QRA� mr 9��#��G��#gWAR�:�BLuq��'4A;88D�A���!I835LD@�PA�A�q3h��!��q3TI���5�β�pgRIA�Q�BAF� P�A���1��5��T����EMJ�I1Q��D�F_�`�ӨQ��LM�t�FA�`HRDY4d�P�`RSoq+`|Q0EMULSE�`x���E� ���I�����$]a-$�Q$�Q�,���� x��EaG�P�AРAAR�2)�09mb�E50��wAXE&�ROB#��W�ac�_�M�SY����Ae�VSWWR�ذ�M12�� STR�"Ņ�d�h�E� !	CUq#��lqBhP3�oV��)��OT�Pv� 	$�ARYg�ЦR_!�`	T�FI���j�$LINK(�1w��Q�_eS3��CU��RXYZ@Q��[��	co��Q�RJ�X�PB!��"Kd0�
 � LcFIeg`3�D�9Ԫ$<�_JN�p"�e��SA�OP_~T2�[53�NqTB�aNB2�bC9��DUQ�BV=6r%TURNb����u�Q�!h�?�gFL�)���B�@+pekZ7�3�I� 1�nPKH�M��BV8r%����c�ORQ&�!�# mX�C�����갦��up��.�<��tOVE�q��Mj�tC�zC��B�W�Fq�� � ��� j�0���qw�P� ���	��q���zC��L5��!ERM��!	v"!E8P���#؄A���id�%"�WP1MP1AX�bP1��&!�Q2� 2!>�\A>���=��`=� p=�ep=��p=��@=� JQ=�@:�@J�@Z� @j�@z�@��@���@��@��ב˙DEBU�$�!�1($�{�P��R�g� � AB�P'N�[��sVְ� 
����Ϥ��Ϥ aڧ$aڧ�aڧqڧ eqڧ�qڧ�A�4�`�2\�RLcLABbb�u� ���1s  ��ER�9P �� $8`� A�!��POB�FЉ�P��ލ�_MRA��� �d O0T<�\�EcRR:�2�0TY��aIA�Vb`,���TOQ+�i�L�@,�7R����� C�A � p�T�P��< _V1ْ.�V�2#cą2\�2k�ȱ��op�8ˠȱu�$W��j6�V�A���$�@"�0,���6�Q�	�@�HELL_CFG��A� 5e Bo_BAS��SR��\p�� �CS�T�1�1��%�22�U32�42�52�62�e72�82��RO ��8��P,`NLzA�cAqB��H �ACK�� >�i���`�`G@���7_PUr�CO�@��OU��P0�W!���3�7LTPX�_KcAR���RE���&@P W1�QUE�� �p9CCST?OPI_AL������PU#�Д���PSE�M���M���T�Y��SO��W�DI�����}�L�1_T}M�MANRQ���PEZV�$KEYSWITCHU#�8��CHE9BE�AT!�E�@LE(�$f�U4�F��5�|K��O_HOM�0�O�#REF�pPR��!)�AUP��C��Op�0ECOư_1`_IOCM�d��������g�@� DH�Q� U۲{�Mw2xQ��p�cFORC�f3 �@��OM�@ � @���3�U[SP�@1��$�@�3�4�14�NPXw_AS�¼ 0��ADD' h�$S�IZ�$VAR\2�D@TIP���
� Ah�аJ�� H�� �BS��AC���%FRIFa��S0e�w	��NF�@�Џ@� x�SI��TEFsj"esSG%L}T�R7p&A�x��#P~STMTJ�2�P�@;VBW�p�SHOW�R��S�V
@�D�� �ԱA005pЁ "� �'� '� '� '5�)6)7)8)9)A)�@'v 'V�	&r`'F(JP�() �P�(,)#`�(F)p�(P`)�p�(z)1�)1�)U1�)1�)1�)1�)U2)2)2)2,)U29)2F)2S)2`)U2m)2z)2�)2�)U2�)2�)2�)2�)U3)3)3)3,)U39)3F)3S)3`)U3m)3z)3�)3�)U3�)3�)3�)3�)U4uI4)4)4,)U49)4F)4S)4`)U4m)4z)4�)4�)U4�)4�)4�)4�)U5uI5)5)5,)U59)5F)5S)5`)U5m)5z)5�)5�)U5�)5�)5�)5�)U6uI6)6)6,)U69)6F)6S)6`)U6m)6z)6�)6�)U6�)6�)6�)6�)U7uI7)7)7,)U79)7F)7S)7`)U7m)7z)7�)7�)U7�)7�)7�)7�$v��VPd�UPD��  ���)�޸�YSLO��� � ���Q���TA�����AcLU�����CUT�z�F��ID_L���HI�IV$F�ILE_�?�+��$��SA��� �hҰk�E_BLC�Kh�x����D_CPU��� ��� �B��T���q�	�R ��G�
PWl�� �LA1S������RUNu�������8�u�?���?�� ��T?�ACC���X -$f�LEN��s���f������I�J�LOW_A�XIh�F1f�,�2���M��	�G�_��Ip��Y�8�թTORn��f��D��ܣ\LACE��Y�f�ٳY��_MA� ��3�	�3�GTCV:�[�	�T� \�{�q�|������	����J����MĴ�JH9�����	�r��2�Ц�������ΠJK�VK��#���#��3�J08�'�JJv/�JJ7�AAL'�P]�/�]�W�4X�5��{�N1����M�I�ڤ�LӠ_��i�a���� `u�GGROU����Bd �NFLIC��R�EQUIRE��E�BU��b�Ŷ��2��c�	�a�� ��� \APPR��C �ܠ
a�EN�\�CLO��l�S_!M`������
a��o� �P MC6�8{�����_MGV�ЁC�l��؎�5���B;RK��NOL����:�R�_LI���$����J��P_�� /��7��{�����6L�O�8��b�>?��� ҍ��z��燡��PATH�������ᒨ��� �$��ͰCN��CA� �]���INe�U�C٠��%�C��UMB.�Y��4��Ez��P���P�7�PAYwLOA�J2L��OR_ANE���L�����������R_F�2LSHRC��L�O��$���2���2�ACRL_�"� �����H�b�$H���CFLEX_����Je�� : r���	�t�����	�������F1����ïկ�����E '�9�K�]�o������� ���$��г�#( ؿ�����TR'�X ˲�`H��% �&�8�J�\�`�i�W�@{ńϖϨϺ���J��� � �����όʁ��AT�ðEMLt �5�J�����JE��CTR,�TN"F�6	�HAND_VB�q_����� $f �F2�֋��SW�^������ $$M���R�ӅH�� �L��E:�FA�������I��A��݀��A��A	��@�۪���UD��D	�P��G	��qYST��yQ��yQN�DY �Z��ּD�E ��)����������H$� � �PT�]�f�o�x����}3>�� {@`��n�vf�ўo�ASYM�������Ͱ����_SH��#�=�'��dLH G�Y�k�}���J��G���gs]y��_VI�/C�x�ӵpV_UCNI���t�#��J� �re�r���t���t� ð	G�(:j��#!PX��A�H��N�3�EB��EN/@��DI	�W#O��iB��N��� � �BI�aAK����吂��U���0`��n�� � -]AME\?0�4g���T��PTpi0��5�����K�,p:��U�I�TKp�� $DUMMY1�!�$PS_RF�� i@$��͑L�A��YPV#��=�?$GLB_T~@���ŕ5���`�CAӁ�c XI�	נ�STȱ��SBR��M2�1_Vɲ8$SV_ER��O��#�SCLߐ�AuO�����0O� � 7D ĐOB���3LO�f�S�y�ÐS��p�1SYSS�ADqR�1��5�TCH�@ � ,f L���oW_NA
�����ă�TSR>��l }J�J ���F��B���G���I ���ID���D���D��� V�p�KYV���bu��� ݻ������);Mt>��XSCREi�W�5�E@�ST��F�#}��a�Ǥ��0u_�0AV�� TI� &����1%������1������O�PISb�1�����UEЄG� �񪠞�SG���1RSM_����U?NEXCEP�����S_ߑ��7��&�p9�T���COU\�ғ� 1֤�U�E��؂6�y�PR�OGM@FL�17$CU&�PO�>���I_�H�� �� 8E��_HE�_������RY ?�0����������OUS �� @��D�$BU�TT/�R����CO�LUM0��s�SE�RV�3��PANE��0V���TpGE�UA|�F��ʡ)$�HELP��bETER5�)��E���Oq ��30��;0��M`��U`���]`��IN��-��TpNp��0�131�� �i�L�N��� �0���_�����$H_�0T�EX�3j�^�~$RELV"D��~Ӑ�jb���Ms�?,���p��4�򪑥#��U�SRVIEWV��S <���U"�]@�NFI�0��FOC�UA���PRI�`�m��h� TRIP>��m�UN��Є�� �`/��WA�RN����SRTO�L��&�Rs�O��cORNsRAU�W�vT�	���VI��υ� $���PATH���CwACHV#LOG��LIM�r�S���BR'HOSTǢ�!���R|�OB�OTƣ#IM� ��Si@�0r��������VCPU_A�VAIL���EX
�!�aN��} ~�Ma0�Ua�]a �����ƀ$BACKLAS� �!�$"W���  ��CT%s��@$TOOLǤ$ޮ_JMP�� y���$SS�|v4iAVSHIF`у�PB���Ǥ���Rk(�OSURz�3W�RADI�$��_���%�м1��ぺ��$LU�q$�OUTPUT_BM��IM���b� �}p���#TIL�'SCO�"�#C���$N �&N�'N6N7N#8���u%=,�2�eb`V��υ�<��DJUrU��P_�WAIT���<���:%0NE~���YBOW� ��� $������S�B"ITPEo�NEC/,B@D(D�PJǐp�Rv hE(�#=@�0�B�E/�M�KT����"y�� An�!�OP��
MAS��_DO*آ�qT��D]�����C��RDELAY��SJO�"X֡ �c'T�3��`� ��,l�y�Y_RI wR�#ƢA�? ޳1ZABC�� ���R��
����$$C�X�����Q�����P�PV�IRT�_�PAB�S�!��1 �U�� < �Q(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�K�|`�AXLMTZvK��c  �]��INf�x�\�PREȏNk�����LA�RMRECOV ��Y�����@F ��U�QdK��"�4�F�T����w���������,��P$o�X�NGu �k	 A  � �,�`PPLIMCu�?�U����Handl�ingTool �m� 
V7.7�0P/36+���
��_SWr�Fy0���� 43�����yϋ�7DA7��철
f��r�m�None����Oհ�P�T����<�_+�V詥R�v�7�UTO�RX l���n�HGA�PON�Pe� an�U�' D 1�� �и�����T�n�� oQ 1�  ��*������	7�H帵�]��R�R g�a�,�H����B�HTTHKYV��R�+�=�O�� ����3����!�?�E� W�i�{����������� /��;ASe w�����+� 7=Oas� ����'/�// 3/9/K/]/o/�/�/�/ �/�/#?�/�/?/?5? G?Y?k?}?�?�?�?�? O�?�?O+O1OCOUO gOyO�O�O�O�O_�O �O	_'_-_?_Q_c_u_ �_�_�_�_o�_�_o #o)o;oMo_oqo�o�o �o�o�o�o% 7I[m��� �����!�[����TO�C�U�DO_CLEAN��5Ի�_NM  	�Կ���+�=�O���_D?SPDRYR��HIa��@����ϟ ����)�;�M�_�pq�������MAX@� ��[����׳�X������҂�7�PLUGGp�У���S�PRCt�B���������O�}�5�SEGF{�KY�k�v�������Ͽ���=�p�LAP����o�Y�k�}Ϗ� �ϳ�����������|1�v�TOTALզ|��v�USENU����� ���ߎ���R�G_STRING� 1s�
�kMl�S3�
�ѿ_ITEM1��  n3������"�4� F�X�j�|��������������0�B��I/O SIG�NAL��Tr�yout Mod�e��Inp��S�imulated���Out���OVERR�� =� 100��In� cycl�����Prog Abo�r����~�Sta�tus��	Hea�rtbeat��MH FaulAler%	U�C Ugy������ ���۞��� �6HZl~�� �����/ /2/�D/V/h/z/�WOR y��۲!&�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO0NPO��V@�+ ?OyO�O�O�O�O�O�O �O	__-_?_Q_c_u_��_�_�_�_�_QBDEVYN�PmO�_!o3oEo Woio{o�o�o�o�o�o �o�o/ASe>wPALT�q �/x����� � 2�D�V�h�z��������ԏ���
��GRI����B���j�|� ������ğ֟���� �0�B�T�f�x�������0�j�R�Z��� � �2�D�V�h�z��� ����¿Կ���
���.�@�R�ԯPREG �~����dϲ������� ����0�B�T�f�x� �ߜ߮���������X���$ARG_� D ?	���9���  �	$X�	[�M�]M��X�n�,�S�BN_CONFIOG 9�������CII_SA_VE  X������,�TCELLSETUP 9��%  OME_I�OX�X�%MOV�_H����REP��S�&�UTOBA�CK�����FRA:\x�c Z�x���'`��qxǣ�l�INI�p�x���l�MESSAG������A�>��ODE_D���ă�#O�P2l�PA�USVA!�9� ((O<��� ����� (^L�p��e~j@TSK  ux����o�UPDT) ���d ?WSMg_CF��8����%�+!GRP 2
V5+ L�B��A��#�XSCRD/!1�5+ ����� ��/�/�/??(?�� ���/p?�?�?�?�?�? 5?�?Y?O$O6OHOZO�lO�?O(�r�GRO�UN S�CUP_kNA�8�	r�n�F_ED��15+�
 �%-BCKEDT-�O0�%_LI_�� ���-r�_x�o�o�x���U2r_/��_�_�R��o�iU�_&o�_�_ED3o�_�o�_n_o8�o9oKoED4�oro�'�onn�o�oED5^�:n�8���ED6���o��nK���%�7�ED7��^����n�8Z�ɏۏED8J�*_��N_m����m���ED9�[�ʟ`m7����#�CR_ ����7�ٯD���ū��@�@NO_DEL��O�BGE_UNU�SE�O�DLAL_?OUT ��R��AWD_ABOR��𦾦AݰITR_�RTN����NO�NSi ����C�AM_PARAM� 19�#
 8�
SONY X�C-56 234�567890H ���@���?}��( АZʨ��yŀ��\�H�R5o�������R5y7����Aff�� \�L�^�Z��ߔ�o߸� �ߥ��� ���$�6���Z�l�a�CE_RIWA_I(%;��F�!{�x� ��_LIS$�c%����@<��F@�G�P 1Ż����OK�]�o�.�Cg*  ����C1��9��@��G���CVP C]��d��l��Es��R������[��Um��v�������_�� C���& ���G��;�HEנO�NFI���@G_�PRI 1Ż ��T�������� �CHKPA�US� 1I� ,�BTfx� ������//�,/>/P/b/t/�/Oƭ����8�!_MkOR��� ��@�B�%���?�;̋��	 �"�/ :�/.?9��;P=45��"����-=ֱ?$99��3�@K�4���<P������a�-8��?OO�J
�?KO�'ưS�P1���:O��i`��PDB� �-+�)
mc�:cpmidbg��Od��C:�  &%#P$���Ep�O-_��C  �0	
0
V�@�Oq_<Z��  ��P�0S[_�_=Y�װ���=S[g�_o�\ �� WS[f�_KoA�Mo�JDEF �ch�)�B:`buf.txtqo�Mro��0����'�	�A�ޙ1=L���jMC
�#�-,���>ss��$�-�r���Cz�  BH3Cs7� C���C�M��F��iDP��E�~�WJ!0D��tE�qaE�pIJ$�3H?HƷ��{�G�G��G�G���N[5�K~w)L��X�WI��>�fu7���4�),�,�.װ��,�,��@�u�K�)x6�q�* �* e�3D�n��pEWL!0�EX�EQ��EJP F�E��F� G���}F^F E��� FB� H,-� Ge��H3Y���z���33 '�T5WDn6�P1�@��5Y���"��A��1WDq<#�
 ��O+�)�Zj�bRS/MOFS���n6���iT1� DE � �?DR 
�,�;�&�  @�:��n/TEST�bo�8�ER��!�/3�nvC+�SA�WJq� [���rq�C�pB1 w�CRy�@T�6��T��FPROG %ź��ů��I������喤KEY_TB�L  �6Q�!� ��	
�� �!"#$%&'(�)*+,-./0�1g�:;<=>?�@ABC�`GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~��������������������������������������������������������������������������������͓���������������������������������耇�������������������s����LCK�xX	���STAT*���_AUTO_D�O���G_�IND�T_ENBK��"R���i�[�T2��\S�TOP���"TRL^��LETE�����_SCREEN �"�kcs�c��U��MMEN�U 1""�  <����|�WE[� �ߺ�V��߽������� ,���b�9�K�q�� ������������� %�^�5�G���k�}��� ����������H 1~Ug���� ���2	Az Qc������ �.///d/;/M/�/ q/�/�/�/�/�/?�/ ?N?%?7?]?�?m?? �?�?�?O�?�?OJO�!O3O�OWi;�_MA�NUAL�Ϟ�DB;CO��RIG�4ɟDBNUM�`��<q*�
�APXWO_RK 1#"�ޟ�+_=_L�^_p_�[�AT;B_�� $"���ipT�A_AWAYz�C
�GCP *�9=���V_AL�@Mτ�R�BY���*��H_�` 1���� , 
^7�6�Boo��f�PM��Ij��\@|��cONTIMכ�*���fi
��$cMOTNEN�D�#dRECOR/D 1+"�er9�Q�O�Oq=6��R {���Hx��O �s(�:�L����� ����ʏ܏� ��� $���H���l�~����� �Ɵ5��Y�� �2� D���h�ן������¯ ԯ�U�
�y����R� d�v����������?� ����*ϙ�N�9�G� �ϧ`�^�ϼ���=��� ����(ߗϩ�^�p��� ������9�K� �� ��!�H��l����ߢ� ��K�a���Y��}���D�V�h���RTOL�ERENC�TB��b�PL���@CS_CFG ,0k��gdMC:\���L%04d.C�SVi��Pc���cA� CH z�P�oo�n"W^m�c��R�C_OUT -�[=`�o��SGN� .�Ur��#��25-MA�Y-20 15:�37 �Q�
1:0�0 af P��X��n �p�a�m��PJ�P�{VERS�ION �
�V2.0.11��kEFLOGIC� 1/�[ 	�tH�P��P��PROG_ENB�_\r�ULS�g �V��_WRSTJ�N�`�Fr�TEMO�_OPT_SL �?	�Uac
 	�R575�cO 7�4T)6U(7U'50y(t"2U$tH�/z>2$TO  >-l�/{V_�`EX�G�du3PATHw A�
A\�/�]?o?�kICT	aF��P00g�Tdc�eg��1ST?BF_TTS�h�I��3U�Cda�6�@M�AU ��bMSW��10i�<�l� ��2�Z!�mO|3bO�O��O�O�O�O�O_tSBL_FAUL� �3�_�cQGPMSyK��bTDIA��4�=�d`��a�1234567G890�Wc|6P�/ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�oh�o\SpPf_ *��OR*�?%�PBh z������� 
��.�@�R�d�v�H|Έ�UMP4!Y )^��TRNBKS��Ā�PME�5ЏY_T�EMP��È�3p��D3����UNI.���YN_BRK �5����EMGDI_STA%�W��NC2_SCR 6G��_����͟ ߟ�f����0�B���~�e�17��;�������¯,R|�d�8G��a�������N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶�0������ @$<��)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� �����������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/��/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgO�/�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo�Oqo �o�o�o�o�o�o�o %7I[m� �������!� [oE�W�i�{������� ÏՏ�����/�A� S�e�w���������ק�ETMODE 1�97�v� �'�� �W�RRO�R_PROG �%�%���X�'�TABLE  ��A�������њRR�SEV_NUM ���  ����)�_AUTO_ENB  #���j�_NO� �:�
��  �*�F��F��F��F���+E�_�q�����HIS�h���_�ALM 1;�� ���F�F�+ �� ��$�6�H�Zψ��_�%�  ��D����ېTCP_�VER !�!�F�j�$EXTLO�G_REQ������SIZ����T�OL  h�Dzި��A ��_B�WD�5��a�	�_�DIO� <7���	�h��k�ST�EPw߉�ې��OP�_DO��4�(�F�ACTORY_T�UN��d��EAT?URE =7�a���Han�dlingToo�l 7� DER �Englis�h Dictio�nary=�7 (�RAA Vi�sS� Masteyr0�>�
TEa��nalog I/yO7�>�p1
a��uto Soft�ware Upd7ate�� "`���matic Ba�ckup;�d
�!��ground Edits��  25L�Camera��Fމ� "Lo��elyl��>�L, P��7ommj�sh�8�oh600%�co�����uct%���pa{ne6� DIFD��'�tyle seolect�- `��Con��j�oni�tor<�B�H��t�r5�Reliab��� �(R-D?iagnos����:�y�Dual C�heck Safety UIF���Enhanced� Rob Ser�v��q (V��User Fr����T_iE�xt�. DIO ��f�i�� Z�\=en]d Err��L��O  pr�[r���C  P���EN�FCTN Men�u��v����.fd�� TP Inp�f�ac�  
v�G���pl�k Exc�	 g5t��Hig�h-Spe Sk}i��  Par\��H��G mmuni�c��ons��\a�pur� p���t�\h8��c�onn��2� !�D�Incr� stqrZ�i�<�M-6< �KAREL Cmod. L� ua����8sRun-T]i4 Env=�(m�qz m�+��s��S�/W=�"y�L?icense��'� a���ogBo�ok(Syo�m)�:��"MAC�ROs,�/Of�fse��f���H�G R��M1?�Me�chStop P�rot��d 5�
$�MieShi�f��9�B6SD�M�ix ���7�y�M�ode Swit�ch��Mo����.J& �M�&��g'� 65�ulti�-T� ����Z�Po=s��Regio��  ! 7Pr�t� Funb>�6isB/1��Num ���dx�P`�312  �Adju:�/23HSM7Z* oY�i8�tatu1<�AD� RDMot�N�scoveW� �#��3�uest 867.�9�oG � �SNPX� b����Z#Li�brV�;�rt IDE,� S$@�.�0��� �s in �VCCM9��0��� ��!9�3��/�I� 710< TMILIB�MJ0,@�� �Acc����C{/2@�TPTX"+QTeln �Lq�3�%|(PCUnexcept /motn�� �0�0�,	7�\m72�f�+4�f�K  �h64aVSP CSXC9�@(P�U["�3� RIN�We�'50,D��Rv9r�	menS@� �QiP^ a0��3�fGrid�1pl?ay F O`�f�p@��vVM-�@A(_B201 f`2�� ORD|�sci�i��load3�4�1%�lJ�i�Gua�r�dP�mP��k7��b]aPat�& 0N"Cyc��0gori���`iC00oData�@qug��c�3[,`�3FR�LOAam�5<�3H_MI De�2(�1noc644�0PC�~sePasswo�aA)qp�1p���{-+PvenjCT����YELLOW B�O�I t�"ArcV0vis���%����Weld� cia}l�$    �e�t�OpA ;�41Y\\�5a 2��a���po)@`@�aT14���50.2HT� @ 3xy�R:�82��`g�P��xp�� 1�2�AJPN ARCPSU PR\A��TEh0OLwpS;upg�fil5p�Qp��^ l�cro�6 "T�`�3ELdx�!��SSwpeet�ex^$ J3�QS�o�t� ssag&�% T�eBP� ] <!9M�Virt��3�9�V h	`stdp�n6��ro� SH�AD�pMOVE �TF MOS O �� Dget_�var fail3s ��ߐ  � D���E��� Hol�d BustdCV�IS UPDAT�E IR��CHM�A 62�q�WE�LDT�@S ) �"���: R74�1-�ou
�b��m� BACKGR�OUND EDI{T Ò m41�0�REPTCD C�AN CRASH� FRVRTO�C�ra.�s 2-D���r �0r$�FNO NOT {RE��RED �o PCVl�JO�P� QUICK�O�P FLEN .�pc�c���TI{MQV3 ldm�P?FPLN: 燹 �pl 2���FMD� DEVICE �ASSERT W�IT iC��sA�NġACCESSW M �aŀo1GQui��<!�C"��USBU@- t &? remov��<��2� SMB NUqLApܡ��FIXW�n�HIN͑OL2��MO OPTt�POPOSTwp��D��s- � �Add���ad. 	�io��$�P:�Wu`.$ѠO���IN��M��CP�:fix CPM�O-046 is�sue�tJСO-�|�2�130���S�ET VARIA�BLESΐ�$O�3�D m�"viewc da`PWea��80b. of FD� ��u)��x O�S-1�p� h s� v�D�5t��s Υ�lo �(� W�Ax��"3 CNTg0 T�S$Im��Z#ca��PSPO�T:Wh�p��s�S�TY܄At�pt��do GET_�l���VMGR L]O�0REA�pC��M`P�@ Y��0�_ELECT��L���ING IMPR� N���Rɰ̐sP�ROGRAM�R�IPE:STAR{TU�@AIN-��|D��QASCII�d�OF L���!`PPTTB: N���MLKdme�4��:v�moW�all���R� Nu�Qr� A#ng���`d���tho�n[� ch� >`ܐ�r R2to�un�H85@�iR�CalA�"Sig�n�0�pI,A�Thresh123�#�.c�Hڰ : �MSG_P�єpe�r �ࠡ��A�z�ero5P� A�  �J�!O�Imr � 2�D�0rc imm��`SOME�s�O�N������0SRE�G:�^5� LB� A9�KANJI&H�no��`c	���n dq�� -1�o��INISITALIZATI���we��0= d�r\  f��aP���m�inim90rec� 1lc0�:?!b7lem��ro��L�4<3a i� 09 ��*b�d�w-� ݡ��0�w uHQm@se�4SY�M��s����QЧ 090�WluZ� E;BRe��jձ24�1���m ���P�ar�r@ G�Box fo TME��ːRWRI<���S�Y��\k��F/�u�p��de-rel�a2Qd��#5�bewtwe�pIND���GigE sna�p�us5�spo� V�TPD��D�Os�ġHANDL� �`�Q�i�D��n�0 f.v���B�operabil��` tmCQ��: �H5@�`l��L�
!� ��m@ph�so UIFL�PO>��FA����ΑV7.n��CGT��pi�A�sM�5pj�)@U��i�ne-RemarykO@0 RM-�$�ÔPATH SA̐LOOS���v�`�fig�GLA � �0%���p��J� yki q�ther�An� Tr�`in�D�W����2�7�� X��е���8`n;� IC� ��:  6�d� �y* it 35\�k�Pay�a[2y]_�D1: g��s> dowD2	SD�ISp�1�EMCHK EXCE ֠��$MF +  ��hD�"�P��Վ�B0� ce1Ȣ��me�� �c� !?��b<P�� BUG��yB�
�@DŠPET���V0�0�T93X�X�PANSI)�DI�G��O  H5��P�CCRG E�NCCEMENT�`�Mm�K 1A�H� GUNCHG �OA�1Tڐ����S�g\d���10ORYLEAK�������LC WRDNk R��O�`j5`PNO�SPEްCG��V ont��VM�����W��@`GRI�,@A�7��� �PM�C ETH�0i�SyUذ>� H57�P^0PENS!�N��|��ː RE (i��ROW<�³RMV ADD  II��=p��DC^ q�T3� ALAӀ ��m���VGN EAR#LY>���f n� ��8衸E�ALAY7u��R�PDg�ˀH1SS8�OUCH��D��F�h�����PCDERR�OR*PDE��� W{RO��CURS�P:ٰIp@N gҰ�^?Q-158Kwa��N�SR �ġU3���\aptp��@T�RF@�R�\`�UB��U �`��#RB�0S?Y RUNN���`�10�ఱBRKCT@qROq�Ԁ��ІCDAX��Djj�EISSUcހ\��D��WTSI�aK�tXM��IPSAFETY� CDECK "M6���dѤ�[`S �U�)��4}P@QTWD���E�'QINV��D ZO����a�sb_aBDUAL@|�'QJòF��E�4l�6���P`NDEX F��P�U���SUF�rP�k�Lbѳ�RRVO1/17 Ay�T���ܤ ��FAL�BTP'247���P?q�EwHIG�PCC n���0�ESNPX*PMM�Q ��)!SQ�"�V��8T�bDC�BDE7TEC��ds!Sˀ�BRU/b63���s� 02"�t�s�'�!Ih� Z�T�7pS��"e���߆��,����߉ـ�0�
ա��ق�cscr�ـ �dctrld.؁����fّ��!ĺ��fـ*��87�8��-�% ��� Krm��
�Q�R��78�RIـA�̑ (��~��Q.����ao�ـ\��a:P����a��I��ta 3 "K:����<�#�o���tp؁ "PL�CF"E!�ـ�plcf���ـ-����mai�ـN���ovc���ـt�/�ـ�������􁢐r67�4��Shape GGenwـI��R,���ـT�іV�c (5�ـ��II����� �+��ـl���suga 4P� 4j��I�r6ـŲ5=�5�ѺI���ets6� e" PC���nga�GCREѿ|�5��@�DATj���5ŝ�#t.!��5�a񯜳>A�gtpadb���Y�tput��������ñ��2ـ��5Ę������sl�q� 7�hexy��4�8����2�keyy�ـ�"�pm������us9ߜ�gcـ�����+�H�a�j92�1��pl.ColAly󔱾�r�ВN���ڕr� ({�ـip����r��'���8�7�=�7���tp�� "TCLSj�|���clsk��D���s�kck���)�U�������r�H���71�a�- KAREL Use Sp�POFCTNj��7��a�a��� (��ѡ��@ �ـ��ٹ�6�8=�8"   �ـ� 0S�(V�   lm� 6�99�~ F�)v�mcclmf�CL�Ml��`��60vet����LM:����s�p]��mc_mot���ـy���suX��60���joiT�J��_logH���trc��ve�%�� �����g�f�inder��Ce?nter Fb!��M�520����g��  (m)r,���fi��1��a#z�`� �ـJ��$tq�? "FNDR���~�$etguid@�UID�ـ
?1��pE7�q1nufl��6 �ـ>_z #ѯ7A�x��(�2#<���$fndr����c$��tcpS$]�C�P M� H�3ـ5317��g�38�vC �gD�*Y=�F| Ց`� ^ ���CtmgA4�P��O�CG1ՑO7`�Y��8�Etm �?�Wـe�?�C�Rex�ے���Z����Xprm؁�_�D�_vars�_Z$M ���Vh@����`�gG���ma�w�Grou�p�@sk Exc�hang{@ـÖM�ASK H5�H�593 Ha�H5����`6�`58�a9R�a8�B�a4q2��"�b(�o#
k�/��(�`hp8�0Y0/_��t�qTASKY_�r�$�pz�h�Z�m@���������SDispl/ayIm��v{Gـjʑ8�OJq(P%����@a���a��� ـlqvl "�DQVL�t���q �����Ϧ�y�����1avrdq֏4ᩅ�sim���0��st��o��d���������v�0Z樁���"v��Easy Nor�mal Util�(in4�|+11 J553��a�c���(���0��)�M�<�O��<� k986TA8���#�4�� "NO�R�
��1�_���|�su��.������7����a!g�y! menu�u��g#M�����Rw577� 90 ̒oJ989��49�Lt�A0�(�ity�E��A�,�P�m&��m	h8��"8 2��܄�����C8_Sշ�n? "MHMN�r%. Ը%���ͯ�s����i�Ը-at�Х_����0���ֶ��tm�?м"z�1����Q�2�Ͽ��z�3zos�odst���
�mn�O��e�nsu�Lm���h�RaL�߃��hus�erp�a����c ~���Ը5�ɯ������oper���XԸdetbo`Ý~ �� LUA��������?dspweb����+�X���u<1��10!1W�הּ�2N�A��e�30A#0����4N�;2e�5��|����"��CalxN�0�O ��Z��0�O�$�S%j{��u��� 0Ss�}���ump��\bbk968�!�68�!��b�eq969�9�%��F0�b�� "BBOX��ۍ�schedx����setu~Xk��� ffH)�0��eq)��0�ccol(�1bxc��8�li�Љ�aI����W!i�e@m�rof$TP EB!TA&@ry|M427�*l!s(T\�Q!RecX" H
�qz�?$it%�?#�сk971�!71��{�F�$parecjo��A��?'�����Xrail�@n�age��~@]��D2E� [0 (?:H͒V|x@1ipMa���3�p�!4�"4�u��3�paxrmr "�XRM$��3�rf�Ͼß1�1ꫝ0�y?turbsp'G#8��^@ �015: ��625t/~A��\BH��'ZDiy!:k�E�6@�"A���H� �7���P�.�E!pd "�TSPD�}�T�GtsglD��kY��O�CiCsRct%���HvrvQ���K�P,�~�A  q�#-a21�Y@�AAVM �r-b0� �fdE`TUP� him (J545 l) ��i`616 V2�VCAM .�CLIO Y10uk 5W` (F�`OMSC ���bPs�?STYL�Sua�28 kr�`NRE� I��`SCHgRp�DCSU t�psh ORgSR �ua04��EIOCW`\�fx�`542 L�EX"�`ESET���iay`0shi`7�y`"RMASK��b7o�-`OCO[�x�a7p3Sv q`t�7p0kv6U`xv39�_v�xLCHRvOP�LG�w03;uMHCR3MpC�`YaP`��p6�.fia54�; #�MpDSW�`5�88�ip1�a37� 88 (Dr0�c�5r4���r7 q�j5r5�5r^v�p5��"9PRST� VRFRDM�C�S�a��-`930� ��`NBA  �g1�`HLB 3 �(�aSM�� Co}n�`SPVC L�ia20�#-`TCP� aram\�TMIL r�P�ACC�TPTX ��p�`TELN �96�0�r9/uUE�CK�1r�`UFR�M etL�aOR� ���`IPLKeC�SXC�pj�qCV�VF l F7�H?TTP strbZ0�zcpCGy�8�AIGUI�p7 ���PGS Tool��`H863 dj���qM�Oq3
vJ684c�\$���sPق�s'�1ےs�a96 TFADȑ�651�Cq53 V� oo�b1�44r�-�k�r9�VAT>��J775 �R�=6uAWSMے�`CTOP �q�`�old��a80;!d�iy�XYY�0 ye��i`885 '�B�`L�`u"�`� 7H�`LCMKP��pTSS J%�
�W��CPE \di}s�`FVRC m���NL�U002� 
�en%�6 6i5Jr'�7[�U0�p!o�ࠠK���t� I��4 URI�5�&�U022 nse�~{�3 APFI�`�{�4�2�`-���ailOP��1C�33O��͐tptsD`U0�40g�43�ٲ4x�۰j� "sw%��1`b	�4�C	�5 ڂ�wx�57�eU0�61��S�6ұro�b9�5g�i��68�����!!��7�w�7�Ё�%���"rke%y��3w��4?ǽ���T���8'�089��U09���P��9�:���2 &�l �9�&�l��9B�VrU185�P�M� slA �!3#�}���1q�0�v4�7��108 	�eэphc ��s�)1�q�4+�1����*A�5/�tx�1���Ņ1]pu�Qѡ�t�1������`��3����6���1!p �`�о�-� W8�147 ase C�U`sB�/1 82��1�4~�8 (Wai���59 ��aU16$6�W�1�W�4� j �U�6�#U�7�3U�8 �3ѱ��B��1{���2 act���6 �"MCR@�ِ4�1p������967ǑOU193�3��6��2Y�sP��2A��21��as�F����<�2-���E�2 wDF���55�(��� ��cر5)�w���q��p����qf��L��$� �����q4d��2g�8q��8�51�""]�}�q��< b������B ]�� f�; `�̑� � 8 16 ( ݰ�BA��AAҰ �]���g :�!��>`8 bbfo=�� t� j�� 7 \'� ]�� ��2 k_kv��7�4 &!����W0H5��57&�579s h� L82 %"p��4 3��	5����5��1���594 U219 I7,-�6�p��6i�/\tchH6ur% ��4S3� 90�� h�&�\j670��q���r!�tD�4��&�t6�sg�lc�S�	FrE�H��#F�����hk$��  sC�� ��"F�L�<��dflr��� �� ���fhu!l%�gvPva����sA����"D��3��!creex���!�%�!�%�,����6j6�s�!prs.�!�%�!5��hA�P 5�fsgan��/�/�,at<D��AD���qs`R s�vsch`@Q!Se�rvo S�!ul�eoCA5SVS�!4�4���F��1 (��0Ached�0,`1�EA၍�� �2 Q��0��^�r0�U)1BB�c��� %P5)Q1��V-#�3�1css "ACS�WVY8 8"gA�`8!�/�0��@�e�Ҿ#M��C�3�t�orchm�0�- TQMa�1�1M%�'�9 J5lA59�8 א1�!7)P8 <P(1̢A�ء%R1Qte,�!)E A5E8`ASv�� mLC6wARC_� 1��4q� �V�Ht!tc�A耥Q�4���R F1 7T!2�SEPBPQf-!�RgtmkQ!p@60X��/�PRC8S�Q#�S0�) P�2a96xAn`X�D.<bH5�1�U�}E� T�Qf#` aQ!@<���F!�T!!�a4�3FcRO�Ttm�R!av``58�_�WP��MA$q�E8��>rp�in_����o�@e`Ac�B�rr�)u�!�U�e�td�ѧ�U�Qov�eto�#$,�S�m?monitr42�=�Q�c�st,"M_v�a�P47M��V�0�!� 5�q���ameQ!Ɂrol�A��43$Q0  Sp��16�01$P25�AKR�  �� 0S?�(V�Ɂ)x?j818\nl`mD��zN��r�MPT�P"�O��qmocol�]/
�Y1�4Xa`�@��2�0i�53(1���Touch�!s0ؠ�2%qD2J5 !IU@�٠��= b�0n�� A��]�vP���z�EOLWJ�th��Kwcx���{�etth8!�THSRXâm�t��o "PGIO�sRd�'z�wk� "cWK1�aL&MH�PWH54�5�Q5�o"��m`A��q@7z@6���18�a�PMor��tsn�@T�A�o�c@���"�����m�AuA��T��p�@��T?�|�m4�TM�!2�54�>����m9��w�f��S�3G�qo1r�3���"641��@�8ⱐQ!A�,H E!pRU <�m�Re��h-g "SVGN�_��(copy "COTA��U(��r#j0 "FSG��_�e�h��f�@wA�S�WwjRbY=sgat�u���!�;B�tpN�ATPD7��9 a�79s����sg8!��GAT&o<Rc>9  �Ħ �1�t2`%1�&��1�bpv�1��&�1��B� �1� 6�1�chr`��1�|v�1�sm���1�v���gtdmenps1�(v0!1��mkpdt�r1��]A1��pd��1��$&�1��mvbkup.1��6�A���mkun��G�pr���mkl1�e�P�s1�ni��0&1�l�dvr���glg��t�1��&���#�auth�.p�&��`1�����) sud� 1�7� 1�G�1��\1�g b2�p�w� 1�6O�Ł4�� 1�Ђ   9�46"1����1�t�\paic\p4k9471�wc��|1�ictas-�fMpa�cck0�m	�	gen$!1� wl��Q�9 stfq��q�wb���������vri/�4��^��B1�D��Pfglow�@��Ac0sow�3<R50?�p��Q�TR�  (A0�e T�)B�Ԗ�cu�d!�w�1��z�ac�$046 a� =�f�+paRa���!1�355Ţ1�F�ѡ��)a%��;:afca	ld� �&�0����%�f�m:�"�#�4�`��'a`"�3U���$�B1�! tr�ack���@ain�e/Rail T1rP��{(69�/�@ (L !iEYB�ʔ�_VB!Bu��a 4YB38P�48'7�	�F2��4��/�C�B�1�3Ţ3�/�IUal��1�NT����VA��zQin�p�?0HVaen0�?DXWA�puA�YqBzQtst d�0U�@1GW ��]� j�VD���E&��VH@����openersr^CO�`�ADev/w'~6�F8��񭁶��bA�aes�#1�]� ג�d����m�d�1�k9�@7�6��#�1��/b�epaop`aOPN�Wj�`��Krcel}?�Exg����Y`5Dv��tsc@x?t��a�s Fuvrop /�Dw�nDh��bAr5��QB��g�dk�j!�� Pumpv$Aᛑ�/�1��a;��M��T�q �i���t4U�1�� 0S��O \�mhplug�gr7Gh���u|bZ#��ioh#C{p��v(�AWLIO1�1�@7��S93�Q51�91�t����4�� ST�
yR�t�J989���/RLSE�g1�@C2d�(M�1�/O�'�Q �)�D��G1 zq�H155'?��zq��tcmio��MI�O�$�tc�q"OCL01�UQcP�|�io��u~0%��l9�zp��v�1o����Q�tzt����dtz5I$��V%�rh#�Inte�Q�� C%o~Po�qvRP1�h}d�B554 (l��oBv�,�Q�H��Tcicpc�oo�ڱp5�A�(
��������"Q7`���aڰd�QCD�W�	����8��ڱ�rcnd�_׳1p�a�ײ������S��a��O�2�kz�rpcrt�ᱯ�pٱdEc��S  d�\���u�E!߳vr2k�pE A�-�px�_B\"� choO�l"uC��Y 1খ630@ᗷ�@�� ��`��q��ԑ�GTX�?� �Е1chp "��XOh:�3�&�"85x!E��\p3 � ��P��j�d 11�$h��Plo���҆��ch��3��s 1��a�01���#�Ar��0� !oCB��s�pq[Jm:�k�7�)�vr�Ҿ���a!X%-J�wFRAJ�Watpqrnev'�����fQ��D5�`��KrboT ,�$��PG��[!�sm�ICSP\QQP5y��!QP����j�H[51z�93QP7By�6��������5Ɨ�R6QP���NPR��`(P@aam S�`u�b��ĉa4tpprg�p�B�	�Z�~qratk932(q� v��sc "�iC��~�atp r�_�qqz�;F�LGdsblflt{��ёsable Fau`��CPav��aQ��`aDSB (	Dt$�t�d�A���� QPh"�E1��`f$*��a3[S� A�"tdj � "PaV�Ohf$�1s!bj!��1�"\:1gc���.�f%�du�550�^CAdjust �Point�b��J /��-�0�4�a昐A���j�O�N0\sg��4��w�1\ad=a��"ADJ�M�}j0�etsham��SHAP0���XDjpo �e��G�a��UG�QPG'.��1:�k@ab�5�J�KAR`�ia�gnosti��!<�a��66 J�C��a=P(QL�Q&T�o>�fkrldeP@����	 ��SQ��)�3�/ρ[pp��DBG	2t�!O �U�Rѯ#��V��F( �шS7��Q��ip{�M�ip?per Op��Pq�����78 (MH Gw�1Rlbk_�fTc�BQ��0&�d038�<B8t��E��c�9B_9t��Tc��k����8$q�Sdrnp Vǁ��Qd�Ő6Tea��=���r Mat.Handlv �an`|W�� MPLGv�A_�p�q(�sє�f�� ��g��b��a�� �f������>@$w�� ��Dw��EI d����uu�m���fhn�d "F��  ������#� p��p��>��(Pa�0�To@�$V�!!�3#p�a>��{�Q�k925��26�q�3�{�	p����2	ş�y���7gse>0GS�qďėPR��T���a����tp����{�dm�on_�q�Ŗ�ans���vr��{�=���`��ͪ�<y��wsl�] � pen��D��pY�WA��823X �Q
�G�0!'�&P��8�QqIQ�GQ �\sl��!q��v��� ������֐�_�`����"SEDGiOٳaQ.�tdg�@T�AF8 �F���BN���ÑQm� 7���ڱA��g;Ж��Q�����q�S�ileg�y�e���ϟ�9�F'�QQ�LaQQj517So�3-[JV�?�'�#4A�49GA�W!L�aw {�no�Qf��o�H17D�#a������0t�  �>��LA/NG j�A5��p5�5� gad5��C5�TC5�jp .`5�ce���5�ib=�05��#5���pa5��C�5�WҸ�j539.�f5�]QRu5� Env
5�5S��2K�3y ��J9$5�.� �;��G5�2�D25�JS��p(K>}�n-Tim��"���"��3H􅓹����\kl5�UTIL�"�����r "QMG��,q5�C5��1 "5�ړ5�s5�\kcmn��+����r5���utM�_�l�read���exP����"��\��l$"���135�rt[! -5�tuva��`_�4�5� �`CV�����\p ���Bp9tbox��_q�cycs}kRB�TvveriOPTNv��l���e��K���h�g/�agp.v�1$�"1$ptlit�DPND�BP�m$dn#te\cy�m$8$o"��#mnu!3�/�/�/�.5�/�/�m$��UPDT �ite��.3 sw�to95]�-4oolBD5wb95��-4FR-4Y�� /2grd�-4��-4�b-4��w-4B-4 .3��-4�-4'�-4��.3B0l� /2bx� "�5�Q5I.3t�l�7��AE�#/2r l\�6�@O�-4 :4ColD5eMa-4+�AC�5K�-4W�Q5ml�>-4Chang95}�895�qQ5rcmdE�b�OZ�`6�5,r�7�6¤�7�5&r_+]22�=_O]2� c_u_3U4�<_N^57�_�_1UC�CFM�Ey��_acGcdau59#�6cAE X`�/2|�Da��4|aO/Jm�a�5�-4@ �4�aAOSJ	Q�e�o �oY��-4��ZDQF-4sk��?�@rte�t�q-4\$�3�q�eunc.-4��4�q�5sub�5��5E�q�5cce�@oRf^opm4E�o�fv�7�o�e T �c�o�nt$
Pte;�q �@�f\��k���6;�-4Ѓ �-4K�D��zh!-4xGmov�b�q�et����f�"�tgeo�bdt.���ƥ�e�tu� ɐ��ɐ��t$ɐٓxߟ�z��gvar'��xy&�.�pclJ�cɐ���ɐ�eɐgripssu����uti�|����infpo��ܯ�ɐ�������\����ɐ�Ʊ�8�p���n��ɐ%�ɐZ�m�T���ɐԶ��\�og�ġ�Ʊ�%�p�\�palp�����s����ɐ ݵ��Ŵ����p�p����pkagd�%�7�lclayY�k�A�ɐ��dɐ5�p�������B��|�|�����r��q����rdmͿ���rinT�-�?�s O�Q�c�̿޼s����&��tv�ߧ�h���stn[`��tX01ɐ)�Dɐ� �Tul4�q��g�26Ϥ�upd����#vr����נ1}�3�pנ��ϵ�il3C�FU�l4����T�5e��w�s ߘ�֠�߻�w�cm�(��xfe�rϪ�tlk2pyp��conv��cnvݑ��5�aqg, y�lct���n�p��nit�0���d���(�� � �ɐ 0S��(V�U9a�l �pm�Wse ��2����V�C�� (�z���A�0�|��m����&$��޷'#ro��T/f(&���p1�mI��,��$�+�� �/�)G�?�+�� �L�ɰm ∡P?b6 D�4rg����� ������?�9�� O�7 ������>�/ �T�a�8/�C�����E@��b,֡)?�*��nq?�_9l�-!H���  �HA |��p�QU1 pc! O���P ��S� 	�Q�R@t��`  ?���ɐ8�� �M�.Ore�g.ԃnO�o�99 �� ����$FEAT_INDEX  �S ���P��5`ILECOM�P >���baPa�RUc�SETUP2 �?belb� � N �aUc_AP2BCK 1@bi?  �)�R�o��o  %�o�o�P e`�o)oe�oU�oy ��>�b�	� �-��Q�c����� ����L��p����� ;�ʏ_����$��� H�ݟ�~����7�I� ؟m����� ���ǯV� �z��!���E�ԯi� {�
���.�ÿտd��� ��Ϭ�*�S��w�� �ϭ�<���`���ߖ� +ߺ�O�a��υ�ߩ� 8߶���n���'�9� ��]��߁��"��F� ����|����5���B� k���������T��� x���C��gy �,�P��qi��`P�o 2�`�*.VR�H� *Kq�w��2�PC��� FR6:���/�T@`@/R/�=/|,C`x/�/�*.F5D�/�	��/ <�/<$?�+STM D2M?�X.�E?�=� i�Pendant �Panel�?�+H z?�?j7�?�??-O�*GIF7OaOl5MO
O8O�O�*JPG�O�O�l5�O�O�O5_�
A�RGNAME.D)T?_�o0\S__� �T�_@_	PA�NEL1�_�_%@o0�_o�?�?�_2o�rog`oo/o�o�Z3 �o�og�o�o�oH�Z4zgh%7��KUTPEINS.gXML�o_:\����qCustom� Toolbar�(��PASSW�ORD��FR�S:\k�*� %�Password Config�� ������+��O�ޏ s������8�͟ߟn� ���'���ȟ]�쟁� �z���F�ۯj���� ��5�įY�k������ ��B�T��x�Ϝ�� C�ҿg����ϝ�,��� P����φ�ߪ�?��� ��u�ߙ�(ߒ���^� �߂��)��M���q� ����6���Z�l�� ��%����[����� ����D���h����� 3��W������ @��v�/A �e���*�N �r�/�=/�6/ s//�/&/�/�/\/�/ �/?'?�/K?�/o?�/ ?�?4?�?X?�?�?�? #O�?GOYO�?}OO�O �OBO�OfO�O�O�O1_ �OU_�ON_�__�_>_ �_�_t_	o�_-o?o�_ co�_�oo(o�oLo�o po�o�o;�o_q  �$��Z�~ ���I��m��f� ��2�ǏV������!� ��E�W��{�
���.� @�՟d������/��� S��w������<�ѯ��Ơ�$FILE�_DGBCK 1�@��ʠ��� ( ��)
SUMMAR�Y.DG篓�M�D:�[���D�iag Summ�ary\�i�
CONSLOGQ�4�F����߿n�Console log��h�G�MEMCH�ECKտ��J�c���Memory �Datad�l�� �{)O�HADO�WY�>�P���t�S�hadow Ch�anges��£-���)	FTP�ҿ?���C�n���m�ment TBD�l�l�0<�)ETHERNETa����"�����n�Ethernet ���figurati�on��s�V�DCSVRF`�F�X�q�t��%6� verify allt��£1p�1�DI�FFi�O�a���u�{%��diff����"�6�1������{�� �����	9�CHGDE�W�i����u��&��9�2p������� �����GDM_q�u�.9FY3p���� ���GDUgy/�u�6/�UP?DATES.U ;/~��FRS:\S/��-o�Updates List�/���PSRBWLD'.CM�/��"�/��/��PS_ROBOWEL��g�\?n? ���?���?�?W?�?{? O�?	OFO�?jO�?{O �O/O�OSO�O�O�O_ �OB_T_�Ox__�_+_ �_�_a_�_�_o,o�_ Po�_to�oo�o9o�o �ooo�o(�o!^ �o���G�k  ���6��Z�l�� �����C����y�� ���D�ӏh������� -�Q��������� @�ϟ9�v����)��� Я_������*���N� ݯr������7�̿[� ſϑ�&ϵ�7�\�� ��Ϥ϶�E���i��� ߟ�4���X���Qߎ� ߲�A�����w��� 0�B���f��ߊ��+� ��O���s������>����O�t�������$�FILE_ PRގ ����������MDONLY 1@��~�� 
 �5� Y�0}�=f/�� ��O�s �>�bt�' �K���/�:/ L/�p/��/�/5/�/ Y/�/ ?�/$?�/H?�/ U?~??�?1?�?�?g? �?�? O2O�?VO�?zO �OO�O?O�OcO�O
_~��VISBCK��|����*.VD_|[_�@FR:\F_��^�@Visi�on VD file�_�O�_�_�Oo �O)o�_:o_o�_�oo �o�oHo�olo�o�o 7�o[m(� � D��z��3�E� �i�����.�ÏR� ��������A�ЏR� w����*���џ`�����������O���MR_GRP 1A���L4�C4  ;B�9�	 ��������*u����RHB ���2 ��� �?�� ���ݥ�� �������ި%�ߤA��5���_�J�K���cI��H���IT�RӦ�Q%�'M���q�� Fw'�H>�q�F�p�;����;,� @{����@�iC���iC��E�� Fw@ %5U1����J��NJk��H9�Hu���F!��IP��s��?@�u�ÿ9��<9�8�96C'6<�,6\b���B���$CrC���C2�&B���C&�����A�g�B�	�B|EDA�v��B,fB<��`�������9�A�?� M��r�ߖ߁ߺߥ��O���AG�q@5��߯���� 4��X�C�h��y��`���������BH9�� ��������xC$���F�X�5�
��P�X�P�~����z����ͤ����M�O@�33������\��UUU!U<��	>u.�?!���k�����=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!��7�:�7p��D��@ D�� CY�@�UC���Ώ� ����������/� B/�"/x/�/X�/�/ �/�/�/?�//??S? >?w?b?�?�?�?�?�? �?�?OO=O(OaOsO ��N�P�^O�OZO�O�O _�O+__(_a_L_�_ p_�_�_�_�_�_o�_ 'ooKoXi�Xo~o�o �oi��o�o=o�o�o BT;xc�� �������>� )�b�M���q������� ��ˏ���7�/{/ %/7/��[/��/ܟ��  ��$��H�3�X�~� i�����Ư���կ� ���D�/�h�S���w� �����O㿩�
ϥ�.� �R�=�v�a�sϬϗ� �ϻ�������(�N� 9�r�]ߖ�]o������ �߷o�{�$�J�5�n� U��y��������� ���4��D�j�U��� y��������������� 0T�-��Q�� u������ϟ5G P;t_���� ���//:/%/^/ I/�/m//�/�/�/�/  ?ǿ!?�?Z?E?~? i?�?�?�?�?�?�?�?  OODO/OhOSO�OwO �O�O�O�O��
__._ @_�d_�O�_s_�_�_ �_�_�_o�_o<o'o `oKo�ooo�o�o�o�o �o�o&J5n Yk�k}��� ��1��U���� y���ď���ӏ��� 0��@�f�Q���u��� ��ҟ������,�� P�?q�;?��[���ί ���ݯ��:�%�^� I�[��������ܿǿ  ���6��OZ�l�~� E_Oϴ��������� ��2��V�A�z�e�w� �ߛ��߿������� ,�R�=�v�a���� �������'�I�K� �7�9�?���o����� ������8#\G �k������ �"F1jUg �g������/� /B/-/f/Q/�/u/�/ �/�/�/�/?�/,?? P?;?t?�?MϪ?�?�? ���?Ok?(OOLO3O \O�OiO�O�O�O�O�O �O�O$__H_3_l_W_ �_{_�_�_�_�_�_o �_2oDo�eo/����o e��o���o��
%o. R=vas�� ������(�N� 9�r�]���������ޏ ɏ��׏8�ӏ\�G� ��k�������ڟş�� �"��F�1�C�|�g� ����į�?ԯ���� �?B���;�x�c����� ��ҿ�������>� )�b�M�_Ϙσϼϧ� ��������:�%�^� I߂�Io[o��o�ߣo �o��o3��oZ�u�~� i������������  ��D�/�h�S���w� ����������
��. ����'�s�� ����*N 9r]����� ��/ۯ8/J/\/n/ 5��/��/�/�/�/�/ ?�/ ?F?1?j?U?�? y?�?�?�?�?�?O�? 0OOTO?OxOcO�O�O��O�O���$FNO ����A��
F�0Q P T�1 �D|���@RM_�CHKTYP  ��@����@���@�QOMP_MsIN"P����NP��  X�@SS�B_CFG B��E ���{_��rS�_�_�ET�P_DEF_OW�  ��-R�XI�RCOM!P�_�$�GENOVRD_�DOCV���lT[HRCV deddo_ENB�_ `�RAVC_GRP� 1CdW�Q X �O�o�O�o�o�o�o�o &J1nUg �������"� 	�F�X�?�|�c����� ��֏������0�b�ROUp`I�HQP������R��8�?T쀟3�|��������  D�ڟl���@@�B�������o�4�g`S+MTmcJtm蕗�������AHOSTC�]R1KO�pP��a� M������0�  27�.0G�10�  e'�t���������b��ۿ����4�˿ų	�anonymous8�f�xϊϜϨ����л���%�'��[� 0�B�T�f�x�ǿ�߮� �����Ϗ�E��,�>� P�b������������ �����(�:���^� p��������������  $s����� �������K�  2DVh����� ����5GYk m7/�v/�/�/�/�/ �/�/??*?M/� �r?�?�?�?�	// -/OA?c/8OJO\OnO �O�/�O�O�O�O�OO M?_?4_F_X_j_�?_ �?�?�__%O�_oo 0oBo�Ofoxo�o�o�o �__!_�o,> �_�_�_��o��_� ���So(�:�L�^� p����o��ʏ܏�� �u�١ENT 1=LO� P!��E�  A�3�p�_� ��W���{�ܟ���ß �6���Z��~�A��� e�Ư�������� �� D��h�+�=���a�¿ ��濩�
�Ϳ�@�/� d�'ψ�KϬ�oϸϓ� �����*���N��r� 5ߖ�Y�k��ߏ��߳�����QUICCA0!����p�3�1q�M�_���3�2������!ROUTE�R�����`�!P�CJOGa�<�!�192.168�.0.10:��N�AME !"�!?ROBOT����S_CFG 1K�"� ��Auto-sta�rted`tFTPkH���s� �����$� '9\J���� ��Jv!3E/Y {1/b/t/�/�/g�/ �/�/�/?'/�/:?L? ^?p?�?�?Qcu�? ? OO/$O6OHOZO)? ~O�O�O�O�O�?kO�O _ _2_D_V_�?�?�? �_�O�_O�_�_
oo �O�_Rodovo�o�_�o ?o�o�o�og_y_ �_1�o��_��� ���o�&�8�J�m n��������ȏڏ) ;M_a�F��j�|� ��������֟���� /�ɟßT�f�x����� ����!�#��W�,� >�P�b�t�C������� ο�����(�:�L� ^ϭ���ѯ����� �� ��$�6��Z�l� ~ߐߢ���G��������� ���T_ERR� M��.�>�PDUSIZ   �^���U�>n�W�RD ?����  guest\��������������SCDMN�GRP 2N;X����p���\�KM� 	P01.14 8���   y���}�B    �;���� ����������������������~��\��������|��� � i  � � 
���ҕ������+��������
���l��.V؋�"��luop 
dy��������&�_GROU8�O.M� �	0�p��07�	QUPD � ��U��!T�Y�M�@�TT�P_AUTH 1�PM� <!i?Pendan�������!KAREL:*����KC�����VISION SCET� ://��� Q/?/i/��/{/�/�/��/�/�/"?�/>YC?TRL QM�P��v5��
��FF�F9E3.?��F�RS:DEFAU�LT�<FAN�UC Web S_erver�:
Y ���A<OO*O<ONO�`O<�WR_CON�FIG R<� ��?>�IDL_�CPU_PC�0��Bȩ��@�BH��EMIN�L���DGNR_IOG�|���S�@NPT_SI�M_DOV[T�PMODNTOL�V 3]_PRTY�)X�B�DOLNK 1SM����_�_�_��_�_�_o|RMAS�TEP&|R_O_gCFG"o4iUOD|Eo6bCYCLEdo�4d�0_ASG 19T<���
 o�o �o�o�o!3EW�i{���k�bN�UM{�Q��08`I�PCH�o58`RTRY_CN�0
RQ�6bSCRN>{�Q��U� 6ba`?bU�M��p����$J2�3_DSP_EN� M�ᆀOBP�ROC��LUMiJO�G�1V�@Q�8�?��{}?ŃPOSRE��~VKANJI_` d�
_H��V�W�L}6�h�1�C�CL_L��@�r�H�EYLO�GGINB`����Q�PLANGUA�GE �6�B��4 �>�LGW�X�f?�ҧ���x% �Ԛ�?��@���'0���`$�>MC�:\RSCH\0�0\�?�N_DISP YM�Ĩ�8|�z�<�LOCGR�B�Dz�DA�OGB?OOK Z�kR�`P�T�X���B�T�f�x�����������v6	�<�������_BUF/F 1[�]� I�2��H�S�h�d�n��� �Ͽ϶���������+� "�4�a�X�j�|ߎ߻������ߔ�ˀDCS� ]� =��;���C��5Y�k�}�|���IO 1^�kG t��� ��� ������� �2�D�X� h�z������������� ��
0@Rdxz��EPTM  GdR2���� 0BTfx��� ����//,/>/�)Ĩ SEV:���.�TYP���/0�/�/ �-�RS�0��|*�2�FL 1_��@��9�9?K?]?o?0�?�?�?�/TPѐ���"ݭNGNA�M��p�tU�UPSF��GI���E�A�_LOAD��G [%��%	=AR�0�1�?�JMAXUALRM�w��x{@A�dQ:�<��C��y@C��`��Oj�lM�@̀�Ҁa�k �X�	V�!�p+e���O Τ,RX_C_U_�_7�|_ �_�_�_�_�_oo;o &o_oqoTo�o�o�o�o �o�o�o�o7I, mX�t���� ��!��E�0�i�L� ^�����Ï�����܏ ��A�$�6�w�b��� ����џ��������� �O�:�s�^������� ͯ���ԯ�'��K� 6�o���d�����ɿ�G�D_LDXDIS�A�0���MEMO�_AP�0E ?a+
 � ѹ%� 7�I�[�m�ϑϣ�y@�ISC 1ba+ �����'T,���
� ��C�.�g�Nߋߝ�� �߀�����	���?� ��N�"������ ��b������;�&�_� F��������x����� ��7��F �|���Z�� �3W>{���p���/��_MSTR ca-~%SCD 1d���m/��/|/�/�/ �/�/�/?�/3??W? B?{?f?�?�?�?�?�? �?�?OOAO,O>OwO bO�O�O�O�O�O�O�O __=_(_a_L_�_p_ �_�_�_�_�_o�_'o oKo6o[o�olo�o�o �o�o�o�o�oG 2kV�z��� ����1��U�@��y�/MKCFG �e--��<"LT�ARM_��f�;�� v���|���METPU��n���5)NDS?P_CMNT���8��#�&  g-.a��v���y���#�PO�SCF/�:�PR�PM.� �PSTOoL 1h��4@��<#�
��t���� �����/�q�S�e� ������ݯ��ѯ�����I�+�=��i�#�S�ING_CHK � ǟ$MODA�QӃi��a�����D�EV 	K*	�MC:�HSIZ�E�--ȹ�TAS�K %K*%$1�23456789� V�hŷ�TRIGw 1jK+ lK%3%�a���  ������M#8�YP#���5$���EM_INF� 1kڇ �`)AT&�FV0E0��a�)�I�E0V1&A�3&B1&D2&�S0&C1S0=>P�)ATZaߵ���H����p���	��A�9���]�D��� G߸�k�}ߏߡ�� ��6�m�Z�l���K� ����������� �� ����hs�-����� }����@R v);M_�� �+/*/�N/	/r/ �/k/�/[m�/�� �&?8?�\?�/�?;? E/�?q?�?�?�?O�/ 4O�/�/??�OA?�O �O�?�O�?_�O_B_�)_f_��ONITO�RJ�G ?��  � 	EXEC�1p��R2�X3�X4��X5�Xy��V7�X8
�X9p��R0Bd�R d�Rd�Rd�Rd�R d�Rd�Rdbdb�c2h2'h23h2�?h2Kh2Wh2ch2�oh2{h2�h3h3�'h3�R��R_GR?P_SV 1��>����(q�� �>�EeS�<G����X�����>gc.w�@�_DR�&Λ�PL_NAM�E !��p��!Defaul�t Person�ality (f�rom FD) RR2-q 1m�)deX)dh��q7�X dv� �� $�6�H�Z�l�~����� ��Ə؏���� �2�D�V�h�t�2����� ��Ο�����(�:���<��d�v������� ��Я�����*�踝R,r 1r�yհ=\��, ������f� @D�  &z�?���f�?������A'�6z�ܿ���;�	l��	 ��xJ�԰�����˰ �< ���� ��IpK��K ��K=*��J���J���JV尻�"�ɱT���:�L�Ip@j��@T;fb��f��n���%�4��=�N����I���g��a������*��*  ´�  ��P�>��������n�?z����n���Jm���� 
�ғ�`%��Ī�9��� �`��  P}pQ�}p�}p|  ��r�/׈�+�	'� �� ��I� �  ��J��:�È��È=G�����6Ç�	����I  �n @
�+�l�$��l�!��9�A�7�N�p|�  '��_���@2��@���f�Z��@��C��C�p_C�@ C��C���C��o�
�A��q� "  U@���
0ǉB�p*�A��2���0`�o�R�n�Dz��q���߁�������2���( �� -����������o�' ���!�o�M�� �?�ff ��/A�� ���v�7�a��
>N��  P��2�(o� �e�����ڳڴD�/?��o�x"Ip�<
6b<߈�;܍�<�ê�<� <�&�KNA둳��n�O�?fff?�?y&�3�@�.��J<?�`� M����.ɂ���� �lƴa2//V/A/ z/e/�/�/�/�/�/�/8�F�p�/4?�/�X?�y?�K?�?��E��� E��G+� F���?�?�?�O'OOKO6OoO.�BL��B�_0���O UO[��OcO_o?5_�?�\_�O�_�_�_�_U
��h��V�W>�r_on_/oo,oeoF�GA��d;���CRop�oNoD������o��o%5yķD��f8C|�spCH5�"Z�d����a�q@I��~N'�3A��A�AR1AO��^?�$�?���;��±
=���>����3�?W
=�#���{�e��n�@������{����<���~(�B��u��=B0�������	���H�F�G����G��H��U`E���C��+���I#�I���HD�F���E��RC��j=z�
I���@H�!H��( E<YD09ڏ�׏��� 4��X�C�|�g�y��� ��֟������	�B� T�?�x�c��������� �ϯ���>�)�b� M���q��������˿ ��(��L�7�Iς� mϦϑ��ϵ������ $��H�3�l�Wߐ�{� �ߟ߱��������2� �V�A�z��w��� ����������R�:�q(�q���������e��xv����a3�8���<���a4Mgs�������IB+���a?���{�&&	�fT�x���eP�P��A�O	\�`��*<��R^�p�����  ����*//N/</ r/�)�O� ��/�/�%�Q�/�/�/??'?9?  N?l/�?��?�?�?�?�2 wF�$�Gb��A��@a�`rqC���C@�oTO�dq�|KF�� Dz@��� F�P D��eO�O�I�cO�O�O�__1_�c?��ͫ@@8Z^4� �� �� �n
 8_�_�_�_�_�_�_ oo+o=oOoaoso�o��zuQ ������1��$MSKCFMAP  R5� `6�uQqQ�n�cONREoL  ��a�� �bEXCFEN�Bw
�c�e qFN�C'tJOGOV�LIMwdprd��bKEYwsu��bRUNc|su��bSFSPDTY��p)vu�cSIGN|tT1MOTe�q�b_CE_G�RP 1sR5�c\:�I�2�m���D i���a�Ώ��Ï��� (�ߏ�^������K� ��o�ܟ��ɟ� H���l�~�e���Y�Ư�د�����F�`TCO�M_CFG 1tB�m�V8�J�\�
�__ARC_$r��2yUAP_CPL���6tNOCHEC�K ?�k �׸տ����� /�A�S�e�wωϛϭ��������kNO_WAIT_L�w�e��NT �u�kw[�5�_ERR!�2v�i�� ߠ߄�߾��c���ߴ�T�_MOc�wj�, ���3���PA�RAMd�x�k��tV#���=?�� �=@345678901��������� ���+�U�g�C�����y�������t����UM_RSPA�CE�olV>H�$?ODRDSP��v�2xOFFSET_�CART��yDI�S�yPEN_FILE� jq^�+�v��OPTION_I�O�YPWORK� y'�5s  x�fRuQ��2��2	 �	2���[ RG_DSBOL  R5sx\��zRIENTT5Op!C�oP�a�.A[ UT_SIM�_D��b�b[ V~_ LCT z?��*+^�)�_PEsXE�,&RAT8 �jv2u�p0"� UP S{.�PS0��/��/�/�/�)�$O�2� �m)deX)d�h��X d ��?-???Q?c?u?�? �?�?�?�?�?�?OO�)O;OMO_OqO�O�H2 
?�O�O�O�O�O__1_C_U_%�<�O_�_ �_�_�_�_�_�_o!o�3oEo�O� �Ov 1�r(���(���07�, ��lp�` @D��  �a?��c�a?m�a%�D�c�a����l;�	l�b	 ��x�J�`�o�u��` �< �	p�� �r��H(���H3k7HSM�5G�22G���Gp
������c�Yk|��CR�	>��qȋs�a�����*  ���4�p�p��pT����B_����=j%��t�q� )�/��aD�����~�6  ���UP� Q� �� |�Б�������	'�� � ͂I�� �  ��i�=���������a	���I  �n @)��m�C���m��[��N���  '� ��~q:�pC�C�@�s�p�C���ҟ 5�
���=x@#�7~H9�^�n�B�I�A��Q��� 0�q��bz比������ȯ�����( �� -݂*�΁6���Am� �0rx���m�lp �?�fAfU ܫN�`�����n�8m྿̺>N�  P�aզ(m� ������ q�c�d#/?��m�xA�n��<
6b<߈�;܍�<�ê�<� <�&1j�m�A0��c��ƾn�?fff?0�?y&����@�.���J<?�`�� l�����dѩ�e�ϟg ߋ��d��Q�<�u�`� �߄߽ߨ�������� )� �M�8�q���
���j���f�E�� E��0�G+� F� ������ �F�1�j��U���y�[bB��A ��|����t�z��� 3��T��{����x��t��h��u�w�>��*�`N9K���A��Z�_�Cq�mc��?��//D///
T)���pٞ�a�`#CHT/A
$� !��!@Iܝ�'��3A�A�AR�1AO�^?�$��?�����±�
=ç>�����3�W
=�#��>��+e�� �������{�����<��.(��B�u��=�B0�������	3�\*H�F��G���G���H�U`E����C�+�Y-I#��I��HD��F��E���RC�j=�>
�I��@H��!H�( E<YD0X/�?O�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_s_^_�_�_�_�_ �_�_o�_ o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV h������� �1�C�.�g�R���v� ����ӏ��Џ	��-� �Q�<�u�`������� ϟ���ޟ��;�&��8�q�\�(�����,�����]��������p!3�8����ӯp!4Mgs8����IB+�+���a���{� E�E���s�����Ϳ��J�Pe�P���(�{�4��I�[�իR}Ϗ��ϳ�������  ���˿I�7� m�[ߑ��H� �������������p"�4�F�X�  mߵ���������2� F�$�Gb	��ϲ����!C���@�s�����~ F� Dz/���� F�P DC�����������,>P�?̯��@@W
}�R���������
 W���� &8J\n�p���*� �������1��$PA�RAM_MENU� ?q���  DEFPULSE��	WAITTM�OUT+RCV�/ SHEL�L_WRK.$CUR_STYL ;G,OPT]�]/�PTBr/l"CB/R?_DECSN � �,�/�/�/
???)? R?M?_?q?�?�?�?�?��?�USE_PR_OG %�%�?\#O�3CCR ���6G_HOST !�!;DxO0JAT�BO�C[OmA�C|�O/K_TIME"ܜB�  �GD�EBUG�@��3G�INP_FLMS�K�O(YT��9_*UP+GAUP \��g[�CH6_'XTYPE
����?�?�_o o#o5o^oYoko}o�o �o�o�o�o�o�o6 1CU~y��� ����	��-�V��Q�c�u���*UWOR�D ?	{]	�RS��	PNS2W�V$ڂJO�!���TE�@�VTRA�CECTL 1|vq�� ��_� ����|4��DT Q}q��c�(�D � _ b� p�Uct�dt�et�ft�Ugt�ht�it�jt�Ukt�lt�mt�nt�Uot�pt�qt�rt����  �� �� ��p��p� �p��p��Pv�� v�T� v�t�t�	t�U
t�t�t�t�Et�t��@v�t�Ut�t�t�t�TV�v�t�t�t�At���v�� v�t�At��v�N�v�!t�E"t�#t�'�v�%t�U&t�'t�(t�)t�U*t�+t�,t�-t�U.t�/t�0t�1t�U2t�3t�4t�5t�U6t�7t�8t�9t�U:t�;t�<t�=t�>t�?t�n v�]�v�� v�� v�Dt�Z v�QFt�Pv�Ht�It�QJt��Pv�Lt�Mt�D� v�Ot��@v�Qt�@VPv��v� v�Ut�UVt�Wt�Xt�Yt�UZt�[t�\t�]t�U^t�_t�`t�at� s���������͟ߟ�(�s,�t,�u,�v,�w�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������l���� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_� ���_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� ��_@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/�L/^/h!�$PGT�RACELEN � g!  ���f �|&_�UP ~��e��!� �!� �|!_CFG ��%�#f!� ���$� �/�/;�"DEFSPD ��,�1�� �| IN~� TRL ��-�f 8�%G1PE__CONFI� ��%���!�$�<LID�#��-~�4GRP 1��7�!�g!A ����&fff!A+�33D�� D]�� CÀ A@6B1�f d�$I&I��1�0� 	 p?�"�+@O ´yC[ODKB|@�A�OmOO�O�O�Of!>�T?�
5�O4_F^0_� =��=#�
K_�_G_�_�_�_�_ �_c_�_&o�_6o\oGo�  Dz�c�of 
 qo�oao�o�o�o�o 0T?xcu������IK
V�7.10beta�1�$  A��E/�ӻ�Ay f ,�?!G�C�/>��+���0T����+�BQ�c�A\i�T�D;�{�p�"�B������Ə؏�T�O'O�2�8��\�G���k� ������ڟş���"� �F�1�V�|�g����� į���ӯ���	�B� -�f��ov���K����� �������>�)�b� M�rϘσϼϧ�����<�=�F@ �� '�۫%Wك�W߉ߛ� �6���������%� �I�4�m�X��|�� ����������3�� W�B�{���x������� ������S~� w�8����� �+O:s^ ������
�<�/ /R�d�v�l/~/�ߥ/ ��������/�#?5?  ?Y?D?}?h?�?�?�? �?�?�?�?O
OCO.O gORO�O�O�O�O�O�O �O	_�O-_?_jc_u_ $_�_�_�_�_�_�_�_ oo;o&o_oJo�ono �o�o��(/�ob/ P/&Xj�/��/�/ �/�/��o��3�E� 0�i�T���x�����Տ ��ҏ���/��S�>� w�b�������џ���� ���+�V_O�a���� p�����ͯ���ܯ� '��K�6�o�Z����o �o�o޿*<n D�rk�}Ϩ��� �φ������
�C�U� @�y�dߝ߈��߬��� ������?�*�c�N� ��r��������� 0���;���_�q�\��� �������������� 7"[F����ο ����(�0^� Wi�Ϧϸ�v�r ��/�///S/e/ P/�/t/�/�/�/�/�/ �/�/+??O?:?s?^? �?�?�?�?�?�?�O 'O�?KO6OoO�OlO�O �O�O�O�O�O_�O_ G_2_k_����_�_ �
ooJCoUo ����oL_�o�o�o �o�o?*cu `������� ��;�&�_�J���n� ����ˏݏO�� 7�"�[�F����|��� ��ٟğ���!��� W��_�_�_�����_�_� o���6b�$PL�ID_KNOW_�M  bd��j�#�SV ��3e=�:e��z�����7��¿������j�vmC�M_GRP 1�P���`d�bd@I�߶B�_�
�_��� ��t��@ǘϾ�^��� �ϮϪ�
�����F�� d�(�Zߠ�^����ߔ� �����*��� �f�$� L��Z�|���������,�>�#�MR'Éb.�Tg��� � ���������������� ����Q+%7�� �������� M'!3��������Y�ST'�1W 1�3e3 �i�;0:o A >/g� </N/`/r/�/�/�/�/ �/�/�/?C?&?8?y? \?n?�?�?�?�?�?	O�'2(.:/j��	<=O.3'O9OKO]O�!#4vO�O�O�O!#5 �O�O�O�O!#6_&_8_J_!#7c_u_�_�_�!#8�_�_�_�_!#M_AD  wd3#�x`$PARNUM  ++�5o"WSCHOj ]e
�gppa�i=��eUPDpo��e�t"_CM�P_$�R`ؠ`'�;�)tER_CHK7u��;�Or4F{�RS|�2�#�_MO�Q`��u_�be_R/ES_G' �+-O ���H�;�l�_��� ����Ə���ݏ����w&@�|�5��u u@R�q�v��s�@���� ���sPП����sbP �.�3��s�PN�m�r���s `�������rV �1�P���b@cX���p�$@cW��(��(�@@cV��4���rTHR_�INR|�Taud�<�MASSI� Z�]�MNH�{�MON�_QUEUE Q�.�bvg��g�bdN.pUrqN��`{ΰ�ENDб��EX1E����`BE��ڿ>˳OPTIO׷�{�ΰPROGRAM7 %��%Ͱ���o̲TASK_I�Qd@�OCFG Ꭾ��o����DATuAe���@�2�N�`�r߄ߒ�<� �������ߖ��!�3�xE�W�
�INFOe��"ݘ������� ������)�;�M�_� q����������������n�z�"� �!���OpDIT ���s�WERF�L��#RGADoJ �b
A��0��?��P��IOORITY��av��MPDSPX��eU����OG$ �_TG� K���ET�OE��1�b _(!AFD�E�p���!tcp|��!ud�>�?!icm��nFXY_���b{���)� *J/\/` ���G/�/k% w/�/�/�/�/�/?�/ 2??V?h?O?�?s?�?z�?*�PORT3��Rc���u�_CARTREP�|bk@SKSTA��^�zSSAV���b
�	2500H8�63(�ς5D1�*b`@�����s�O�O�G	PURGE��B�	�yWF�@DO��$�evW�T�a��:WRUP_DE?LAY �bT�R_HOT{��%�o�_TR_NOR�MAL{�}_�_�VS�EMI�_�_oCaQ�SKIP1��u�Cx 	bO\o\@ Jo�o�o�ojh�u�o�g �o�o	�o?-O u��_���� ���;�)�_�q��� I�������ݏ��Ǐ %��I�[�m�3�}������ǟٟ�ͥ�$R�BTIFR�RCgVTM.+D�	��DCR1c�8l����C�xD�OC�T�?ˋ��?9!w<+��em�6���F���·fy���߿��*�1�eo���o <�
6b<߈;�܍�>u.�?!<�&ǯ ���)�ŰHB�T�f� x���������ҿ��� ���>�)�b�Mφ� qσϼϟ�����5�� (�:�L�^�p߂ߔߦ� �������������6� !�Z�E�~��s���� 	������ �2�D�V� h�z������������� ��
��.RdG ������� *<N`r�o �����/�&/ 	//\/��/�/�/�/ �/�/�/�/?"?4?F? X?C/|?g?�?�?�?�? �?�?�?O0Os/TOfO xO�O�O�O�O�O�O�O __,_OP_;_t___ �_�_�_�_�_�_oGO (o:oLo^opo�o�o�o �o�o�o�o�_�_$ H3lW���� �o�� �2�D�V� h�z�������ΈB��GN_ATC 1��O� AT&FV0E0΋�ATDP/6�/9/2/9��ATAΎ,�AT%G1%B9�60�+++�3�,.�Hc�,B�I�O_TYPE  �����ЏRE�FPOS1 1�>�� x��������?�P���� 6�������V�߯z��� �9�Ǜ2 1�����$��� �ƿ<D�ё3 1�^�p������:�%�^�ܿS4 1����Q��������q�S5 1� �ϚϬ���d�O߈��S6 1��/�A��{�������S7 1���������y�|��0�S8 1�G�Y�k��#��G���SMASK 1����  
����e�XN	O��;�A�����͑?MOTE  ��ʔ���_CFG ������̒PL_RA�NG���q��POW_ER ��^ ���SM_DRYP_RG %��%����dTART ��V�
UME_P�ROs� ʔ_E�XEC_ENB � =���GSPD�� #��4TDB�>PRM_PMT�_m�TQ ����O�BOT_NAME� ���׉O�B_ORD_NU�M ?V���H863  ��t ���!\<�  # w	r*!@�"�D|<���PC_T�IMEOUT6 �x��S232
1��� LT�EACH PEN�DAN_ ����e����Main�tenance �Cons�r���*"��/�KCL/C�� :���/? �No Use�e��/U?�v#NPO�218�����t!CH_L� ����7�	�1�;MA�VAIL�a#����t!PACE1 ;2�ٜ �?% dH�9�eF%�<�>�L8�?H �9 �O�?�O�O_�O(_#W TOfOxO�O8_�O�O�_ �_�__o i��4m T_f_x_�_�_�_�_�o �o�oo .�5;A2@NROdovo�o6 �o�o����4��I�N{3]o��� S������ޏ0�Q�8�f�N{4z������� p����8���M�n�U���N{5������ ͟ߟ���%�4�U�� j���r���N{6��Ư د����� �B�Q�r�@5χϨϏϽ�N{7ѿ �������=�_�n߀��Rߤ��߬���N{8 �� ��$�6���Z�|� ���o���������N{�G ��� t���$
�� C� e#p������������� :hL���2��+��^�!dt Y�k���� �����8o R~q���� ��//=/7I km�/���/�/�/ ??+?=?3/]?W/i/܋/�= `�� @NP�5<�?�/�) A�5�?1OCOI?#J$O VO�O�O�O~O�O�O_ �O�O�O_^_ _2_D_ v_�_�_�_�_�_o$o��_�_
o<o~o@oN<
�O�oN{_MODE�  +��iS E�+��ox?v:_��?'y�z	��o��CWORK_AD��m��q�R  +�����p_INTVAL�`�@�zR_OPT�ION1� u���VAT_GRPw 2�+�]�G(���L�� ԏ揥�
��.�@� ��d�v���O�o���d X�ß����ϟ1�C� U�g�)���������ӯ �{�	��-���c� u���I�����Ͽ�� ϛ��;�M�_�!σ� �ϧϹ�{������� %�7���[�m��Aߏ� �����ߛ����!�3� E�W���{����s� ���������/�A�S� e�w������������ ��+��Oas ���?��� �'9K[�����e�$SCAN�_TIM�a��\���R �(�3�0(�L8z�W�p�p
Wt�Z��2#Nq!�#�Y�:.(/1�#"M"2{$!!d�(~!"�!�r #])�0���/�/�/�r�)�/  �P5�0�2 � 8�?U?g?>1D��j?�?�?�?�? �?�?�?O#O5OGO?Nq�%RO�O�O�[N![q;�o�t�Nqp]M�t��Di�t!c{  � lM"Nq�A !
%�1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�gS�o�o�o '9K]o��� ������#�5� G�Y��o�o�K������ Џ����*�<�N� `�r���������̟ޟ�����1�  0 �B|�_g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ �p���)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� ���ϐ�������� �0�B�T�f�x��� ������������,�0>�P�J�V�  �1�� �������������� 1CUgy��������	 �y3"HZl~ �������C&a5/</+&�r!� 5/q-	12345678R_���L{0�@�/�/�/�/�/?3,?>?P?b?t?�? �?�?�?�?�?'OO (O:OLO^OpO�O�O�O �O�O�?�O __$_6_ H_Z_l_~_�_�_�_�O �_�_�_o o2oDoVo hozo�o�_�o�o�o�o �o
.@Rdv �o������� �*�<�N�`������ ����̏ޏ����&� 8�g�\�n����������ȟڟ����"�+& s�C�U�:�Z���������Cz  Bp�   ���2�/$@��$SCR_�GRP 1�(��e@(�l��� @ >Z! U!m��	  #�-�=�6�n�p�l�S��y(J�w�e������3%Dʰ֠o���ป��M-�10iA 890ƅ%90� Ɓ M61C �#�-I���*#�
\�l�,�O'�|�Z!�S�;�o�}�	�n�����������X �,���Y"N�a� ���ߖ�i�@�.!`/���m�����"��B�BŠ�J�H�a�H�A֠p�  @. ��l��?���D�HŠ����H�F@ F�` �������;�&�K� q�\�������<���`��������B� ��YD}h��� ����
CҾ�?4#��0/v/�%��
��������V��j�@���/ B�*'��P����EL_DEFAU�LT  C�����X!M�IPOWERFL�  P�p%W"} W7FDOe& p%���ERVENT 1O���I�n#=��L!DUM_E�IP��(�j!?AF_INEd ?��!FT�/7>��/[?!K߀? ��J?�?!RPC_OMAIN�?�8��?��?�3VIS�?�9���??O!TP2@P�U6O�)d.O�O!
�PMON_PROXY�O�&ezO�ORB�O�-f�O#_!R�DM_SR��*g_o_!RL(�_�$Yh^_�_!
�0M�O��,i�_o!RL�SYNCo.i8|�_So!ROS�/zl�4Bo�on?�o2S �o�o�o�o5�oY  }D�hz�� ���1�C�
�g�.����R����'ICE_�KL ?%�+ �(%SVCPRG1��������3$�)��4L�Q��5t�y��6����뀁7ğɟ�=��/�9��脆_A��� i������>���� f��끎�	�끶�1� �ޟY������.� ���W�ѿ����� ��!��ϯI����q� �����G����o� ���������9�;� 翹�˂�ҏ䀄��� á������� �9�$� ]�H���~����� ������#��5�Y�D� }�h������������� ��
C.gR� v�����	� -QcN�r� �����/)//�M/��_DEV ��)�MC:�U(��]g$OU�TYB`!x&c(RE�C 1���` � � `  	 *` ` ` ` �!��!U+�#��U/�.D�$`!�"?`!)A�8�+
 �P�b�6 s�'�  �  '� ��    Cf���"�#�!� U` /` �` ��=�y �y �y ���+��` B� D�?O�%��|0��<S  M��H� �0_�k�? O�` ��4)` ��?��T`!y ��0�` k� �NPO�OOc݀;�[0�0�1o  k�=0i�O !� U� �` ` ,` -�xO��y ��!�D�n� M�O]_�Oc��O�@�F��O
__�._@_R_d_If�6r _�H�i@_0�2��x�C�@��_�!er` �\4�P#�_��fy �y �y ��y �` To�ooh}$0k �  � ~�1   �i@�=�o ;@�2�0 l` K`$|o�dy %�y �y Dq��! ,a�oh[�l�0k`��bR  Ȣ l�P
5�2` �` �V(�c�4��D��!ج�ta��; L�  "Ɣ3G�Qݢ �>` �`�� e&` ` w�F���b�D֔DX� >XX��� �aĀ<Đ?g���?�?�?�?���ď"F �;  K#f�4���'�W��  =� �� ��
j` Q� ,���y U�y �H��` U|�b�t��"x1 � �T� B�x�f�������ү�� ����,��P�>�t� ��h�����ο��޿� �(�
�8�^�Lς�p� �ϔ����Ͼ� ���$� �4�Z�H�~�`�rߴ� ���������� �2�� V�D�f�h�z����� ����
���.��R�@� b���j����������� ��*<`N��r�����%V �1��, P 8g@-����*I  W^� e(a*TY�PE�/e"HELL_CFG���&� �q66�0-RS�p ���//?/*/c/ N/�/r/�/�/�/�/�/@?�/)?8;�p:>����` %K?y?�?F=�J1J1�p�>�1�p)��a22!�d�?�?��HK 1�� �a�?AO<ONO`O�O�O �O�O�O�O�O�O__�&_8_a_\_n_�_|OMM ���_FTOV_ENO��nwOW_RE�G_U@�_� IMWAIT�Rq�6k�OUTf iT�IMe��ZoV�AC�1o#a_UNI�T�S�fwMON_�ALIAS ?e~�Y ( he �o�o0��o] o��>���� ��#�5�G�Y�k�� ������ŏ׏����� �1�܏B�g�y����� H���ӟ���	���-� ?�Q�c�u� ������� ϯᯌ���)�;�� _�q�������R�˿ݿ ��Ͼ�7�I�[�m� �*ϣϵ����τ��� �!�3�E���i�{ߍ� �߱�\��������� ��A�S�e�w��4�� ���������+�=� O���s���������f� ����'��K] o�,����� �#5GY} ����p��/ /1/�U/g/y/�/6/ �/�/�/�/�/�/?-? ??Q?c??�?�?�?�? �?z?�?OO)O�?:O _OqO�O�O@O�O�O�O �O_�O%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3o�_Woio{o�o �oJo�o�o�o�o�c��$SMON_D�EFPRO ����4q� *SYS�TEM* . �"vRECALL �?}4y ( ��}!xyzrat�e 11=>de�sktop-b2�5t4o0:10�168 ��q74�4���z}7c�opy md:p�rogram_1�.tp virt:\temp\~@�7�I�[��rsv6} �!���ď֏i�{�� ��0�B�T����� `���ҟ�w�	����� >�P�������+��� ίa�s�������:�L� ^�����'���ʿܿ �����6�H�Z���;��frs:or�derfil.d�at�mpbac�kϏ��������2>��b:*.*�ϛ������8�J�\��6xt�:\��~�ߐ�+�(����a�7t�a|ߎ� ����=�O�b�t����� *������r��� ���P9�K�]��
�� ���#�����������:15916����8 J\o�%�� ����ύ�=O b����*��� r� /�9/K/]/p //&/�/�/�/�  �/5?G?Y?l�~�� �+�?�?�?���ϓ?�( �?8OJO\Oo��O�# +O�O�OaO�߄O�O�  �O=_O_�O�/?_*_ �_�_�_r?�?O(O9o Ko]o�?oo&O�o�o �onO__�O5GY �O�o�_���j/ ��/�1�C�U��z/ ������ӏf���� ����?�Q�d_v_�_� ,���ϟ�t����� ;�M�_��_o�o�o�� ˯ݯpo�����o7�I��[�j��$SNPX�_ASG 1�������� P 0 '�%R[1]@g1.1`���?�j�%��ֿ����ݿ�0� �:�f�Iϊ�m���� ������������P� 3�Z߆�iߪߍߟ��� �������:��/�p� S�z������� � ��
�6��Z�=�O��� s�������������  *V9z]o� ����
��@ #JvY�}�� ��/�*///`/ C/j/�/y/�/�/�/�/ �/�/&?	?J?-???�? c?�?�?�?�?�?�?O �?OFO)OjOMO_O�O �O�O�O�O�O�O�O0_ _:_f_I_�_m__�_ �_�_�_�_o�_oPo 3oZo�oio�o�o�o�o �o�o�o:/p Sz����� � �
�6��Z�=�O��� s���Ə���͏ߏ � �*�V�9�z�]�o��� �����ɟ
����@��#�J�v�Y�r�PAR�AM ����� �	�z�P���j�OFT�_KB_CFG � ����ѤPIN_SIM  ��Ʀ�)�;�ɠr�R�VQSTP_DS�B �Ƣw�����S�R ��� &� ������ΦT�OP_ON_ER/R  ���᱿PTN ���AݲRI�NG_PRM� ���VDT_GR�P 1����  	ʧ��\�nπϒ� �϶���������%�"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�w� t��������������� =:L^p� �����  $6HZl~�� �����/ /2/ D/V/h/�/�/�/�/�/ �/�/�/
??.?U?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFomojo|o�o�o�o �o�o�o�o30ѣ�VPRG_COUNT����^r'ENB)�YuM�s���_UPD 1�>�8  
G�� ���'�"�4�F�o� j�|�������ď֏�� ����G�B�T�f��� ������ןҟ���� �,�>�g�b�t����� ����ί�����?� :�L�^���������Ͽ ʿܿ���$�6�_� Z�l�~ϧϢϴ��������VuYSDEBU)Ghp�p���d�y�SP_PASShu�B?.�LOG [��u�s��9���  ��q��?
MC:\Z�
�[�_MPC`��u��$���q��� �q�ֿSAV �c�؀ԛ�����SV��TEM_TIM�E 1��{ (��p��t�����T1SVGUNS�p�iu'�u���AS�K_OPTION�hp�u�q�q��BC?CFG ��{I�� B��5�` 5�;zC�l�W�i����� ����������2D /hS�w��� ��
�.R= va������ ��/��B/-/f/ Q/�/�/�� �/�/ �/�/�/ ??D?2?T? V?h?�?�?�?�?�?�? 
O�?O@O.OdORO�O vO�O�O�O�O�O_�H �_,_J_\_n_�O�_ �_�_�_�_�_�_o�_ 4o"oXoFo|ojo�o�o �o�o�o�o�oB 0Rxf���� �����>�,�b� _z�������ΏL�� ���(��L�^�p�>� ��������ܟʟ��  �6�$�Z�H�~�l��� ����دƯ��� �� D�2�T�V�h�����¿ x�ڿ�
��.Ϭ�R� @�bψ�vϬϾ��Ϟ� ������<�*�L�N� `ߖ߄ߺߨ������ ���8�&�\�J��n� �����������"� ؿ:�L�j�|������ ��������0�� TBxf���� ���>,b Pr������ /�//(/^/L/�/ 8��/�/�/�/�/l/?  ?"?H?6?l?~?�?^? �?�?�?�?�?�?OO  OVODOzOhO�O�O�O �O�O�O�O_
_@_._ d_R_t_v_�_�_�_�_ �/�_o*o<oNo�_ro `o�o�o�o�o�o�o�o 8&\Jln �������"� �2�X�F�|�j����� ď��ԏ֏���B� �_Z�l�������,�ҟ�������,��J���$TBCSG_G�RP 2���  �J�� 
 ?�   u���q�����ϯ��˯@��)�;�N�U��\��d, �j�?~J�	 HC��8��>����9�CL  B�m�����z�w�β\)���Y  A���B�;��Bl�=�,��ɐ�Z�,��  DA	�{�F�`�j�Cs���όϦϰ̖���@ J��+�>�Q��.�|߀��d�v��������؈�J�	V3.0�0m�	m61c��	*,�$�I�;�&D�>���J�(���� r�D�s�  #����D���N�JCFG ���f� i��������������7�E��E�k�V� ��z������������� ��1U@yd� ������ ?*cN`��� ���m����/"/ �U/@/e/�/v/�/�/ �/�/�/	??-?�/Q? <?u?`?�?�?J�6��? ��?�?�?*OONO<O rO`O�O�O�O�O�O�O �O__8_&_H_J_\_ �_�_�_�_�_�_�_�_ o4o"oXoFo|o�o�� �o�obo�o�o�o B0fTv��� ~�����>�P� b�t�.���������̏ Ώ����:�(�^�L� ��p�������ܟʟ � �$��4�6�H�~�l� ����Ư���د�� � �o8�J�\����z��� �����Կ
���.�@� R�d�"ψ�vϬϚϼ� ��������<�*�`� N߄�rߨߖ߸ߺ��� ���&��J�8�n�\� ~����������� �� �"�4�j�X���|� ����n���������0 TBxf��� ����,P >t���d�� ��/(//L/:/p/ ^/�/�/�/�/�/�/�/ ? ?6?$?Z?H?j?�? ~?�?�?�?�?�?�?O O OVO��nO�O�O<O �O�O�O�O�O_
_@_ ._d_v_�_�_X_�_�_ �_�_�_o*o<o�_o ro`o�o�o�o�o�o�o �o8&\J� n������� "��F�4�V�|�j��� ��ď������O�$� �O��f�T���x����� ���ҟ��,���� b�P���t�����ί� ������(�^�L� ��p�����ʿ��ڿ � �$��H�6�l�Z�|� ~ϐ��ϴ�������� 2� �B�h�Vߌ��8� ����rߠ�����.�� R�@�v�d������ ���������N�`� r���>����������� �� J8n\ ������� �4"XFhj| ������/0/ ��H/Z/l//�/�/�/ �/�/�/�/??>?P? b?t?2?�?�?�?�?�?��>  @
C �
FO
B�$TB�JOP_GRP �2��5�?  ?�
G6B�=C�DL��0�xJ�@��
D@ �<� ��@�
D �@@UB	 �C��� �Fb  C��VGUAUA>��͘�E�E�I>��@�A��33=�CLް@fff?�@?�ffB�@Q�E-_8Wz�N��O>�nR�\)�O�@�U���;��hCY�@��  @�@UAB�  A�$_�_�S�U?C�  D�A�LwP�RO�z_�Sb���
:���Bl�P��P�D�Q�_So~
AAə�A�hc�ZQDXg�F�=q��e
o�@�p��b��Q�;�AȾ�@ٙ�@L�CD�	x`�`�o�ojo|o>�B�\u�oh�Qt�s�a@33@QV@C��@�`ew<�o>��D�u*��@� p�qP<{�	�Nr�@@�PZv_p� ���&�:�$�2�`� ��l�&���ʏ���� !�����@�Z�D�R������DT�
Fґ�E	�V3.00�Com61c�D*����DA
�� E�o�E��E���E�F���F!�F�8��FT�F�qe\F�NaF����F�^lF����F�:
F��)F��3G��G��G��G,I&��CH`�C�dT�DU�?D���D��DE(!/�E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[
�F���F��M�;'`;Q���8��`F�O����
F��Q��K�2DE�STPARS  ��8O@3CHRe�A�BLE 1�DK$.�
CP�%� ~ �
P�P�P�	GAP�	P�
P�P���
AUP�P�P�|�'RDI��NA���� ¿Կ���`�Oh�z�@�ϖϨϺ��΀�Sf�LC *ʍߟ߱����� ������/�A�S�e� w���������)M e�iߘ�$���1�C� ���%�7�IȀ�
�NUM  �5UNA�@@ ���[���_CFG ������A@6@IM?EBF_TTk���8LCx�5VERY�6�zK5R 1�DKO
 8�
B@2� �0/�  �� ����� 2 DVhz���� �/�
/S/./@/V/Hd/v/u_��b@L�
6@MI_CHA�NA L �#DB'GLVPCL5A�� ETHERADW ?�550�M���/�/N?0F� RO�UT_ !DJ!��4�?q<SNMAS�K*8LC;1255�.�5��?�?2DOOLOFS_DIk���%9ORQCTRL �mK���hM8WO�O�O�O�O�O �O�O
__._@_�|O�N_`_�_a�PE_D�ETAI8-JPON_SVOFF#O��SP_MON ��J�2�YSTRTCHK �DN�g?�RVTCOM�PAT�X53�T�PFPROG %DJ�%	qaRAM_1x7o�\APLAYl���Z_INST_M��0 �l�W�dUS8_WoibLCK�l�kQUICKME� �#ibSCRE@p}-:tps�@ib�a[p`y�"qp_uy���Ti9SR_GR�P 1�DI ؕ�0��z�@��5�#�Y�G��2  ����S��o����܏ǅ ����)��M�;�q� _�������˟���ݟ���7�%�G�m�	1234567�h����b�XZu1��{�
 �}ipn�l/ՠgen.htm�����*�<��R�Panel� setup@�}�6o��������ȿڿ o�e��$�6�H�Z� l�㿐�ϴ������� ��߅ϗ�D�V�h�z� �ߞ��C�9�����
� �.�@��d��߈�� �������Y�k��*� <�N�`�r������� ��������8�� \n����-�n�UALRM�`G {?DK
  � 	L?pc� ������//�6/�SEV  ��h&�ECF�G ��]�&��A��!   Bȣd
 7/�c-5�/�/�/ ??%?7?I?[?m??h�7t!�r��[ �3(ȏ�?B'Imf?wk�P(%*/O`
OCO.O gORO�OvO�O�O�O�O��O	_�O-_�<�d ��=�?;_I_?pHI�ST 1��Y  �(�  ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,��o�_�_oo ��9 �_�]936�_lo ~o�o�o1b�o�o�o�o %�oI[m ��2����� !��E�W�i�{����� ��@�Տ�����/� ��S�e�w����������L��QL������ 1�C�F�g�y������� ��P����	��-�?� ί�u���������Ͽ ^����)�;�M�ܿ qσϕϧϹ���Z�l� ��%�7�I�[���� �ߣߵ�����ğ֟� !�3�E�W�i�lߍ�� ��������v���/� A�S�e�w�������� ��������+=O as����� ��'9K]o ������� ����5/G/Y/k/}/�/ ��/�/�/�/�/?�/ 1?C?U?g?y?�?�?,? �?�?�?�?	OO�??O QOcOuO�O�O(O�O�O �O�O__)_�OM___ q_�_�_�_6_�_�_�_ oo%o/"/[omoo �o�o�o�_�o�o�o !3�o�oi{�� ��R����/� A��e�w��������� N�`�����+�=�O� ޏs���������͟\�����'�9�K�6o���$UI_PAN�EDATA 1�������  	�}]������ȯگ��� )  �$�ᔒ�O�a�s��� �����Ϳ����� '��K�2�oρ�hϥ�������������� Ha$�7�<�N�`� r߄ߖ��Ϻ�-����� ��&�8�J��n�U� ��y���������� "�	�F�-�j�|�c�������������� +=��a�߅� ����F� 9 ]oV�z� ����/�5/G/ ����}/�/�/�/�/�/ */�/n?1?C?U?g? y?�?�/�?�?�?�?�? 	O�?-OOQOcOJO�O nO�O�O�O�OT/f/_ )_;_M___q_�O�_�_ ?�_�_�_oo%o�_ Io0omoofo�o�o�o �o�o�o�o!3W >{�O _�_��� ���pA��_e�w� ��������&����܏ � �=�O�6�s�Z��� ~���͟���؟�'� ��]�o��������� 
�ۯN����#�5�G� Y�k�ү��v�����׿ �п���1�C�*�g� Nϋϝτ���4�F��� 	��-�?�Qߤ�u߇� ���߽��������l� )��M�_�F��j�� �����������7�0�[�����}�l��� ����������)��$ ��Pbt��� �����( L3p�i������ /(�����$�UI_PANEL�INK 1����  ��  ��}12�34567890 Y/k/}/�/�/�/�$�� W/�/�/??+?=?�/ a?s?�?�?�?�?S9S �*�=��U    �?O(O:OLO^O�?\1 O�O�O�O�O�O�O�O _(_:_L_^_p__~_ �_�_�_�_�_�_�_$o 6oHoZolo~oo�o�o �o�o�o�o�o
2D Vhz$���0��
�E0,/A� M�/�p�S�������ʏ ܏�� ��$�6��Z� l�O����<�?����� T!���1�C�U�g� Z3��������ǯٯ� z��!�3�E�W�i��< ��������C��ÿտ ����Ϥs5�G�Y� k�}Ϗϡ�0������� ���߮�C�U�g�y� �ߝ�,���������	� �-��Q�c�u��� ��:���������)� ��M�_�q��������� (�����~���7I ,mb���� ���3ƞ���� ՟w�������� /��,/>/P/b/t/�/ /�/�/�/�/�/?? ������^?p?�?�?�? �??��?�? OO$O6O HO�?lO~O�O�O�O�O UO�O�O_ _2_D_�O h_z_�_�_�_�_�_c_ �_
oo.o@oRo�_vo �o�o�o�o�o_o�o *<N`��� �������� 8�J�-�n���c����� ȏڏI��m"��F� X�j�|��������/֟ �����0���T�f� x�������?/?A?�o ��,�>�P�b��o�� ������ο�o��� (�:�L�^�p����Ϧ� ��������}��$�6� H�Z�l��ϐߢߴ��� �����ߋ� �2�D�V� h�z�	��������� ��g�.���R�d�G� ��k������������� ��<N1r�� ���;��& 8J=�n���� ��i�/"/4/F/ X/ǯٯ믠/�/�/�/ �/�/?�/0?B?T?f? x?�??�?�?�?�?�? O�?,O>OPObOtO�O �O'O�O�O�O�O__ �O:_L_^_p_�_�_#_ �_�_�_�_ oo$o�_ HoZolo~o�o�o��o �og�o�o 2V hK�o���� ����o�/�/�u���$UI_POSTYPE  �%� 	e������QUICKMEN  ��d������RESTORE� 1ݏ%?  ���,�>�b�m]������� ��Οq����(�:� ݟ^�p�������Q��� ůׯI��$�6�H�Z� ��~�������ƿؿ{� ��� �2�D��Q�c� u�翰��������ϛ� �.�@�R�d�߈ߚ� �߾���{υ����s� %�N�`�r���9�� ���������&�8�J� \�n��{�������� ����"��FXj |��C�������SCREր?�ۍu1s]c'�u2G3GU4G5G6G7Gy8G��USER)d.@T(IksQ��4�5�6�7�8���NDO_�CFG ޖ� � &� ��PDA�TE ��None V���SEUFRAME�  ��&!R�TOL_ABRT81/��H#ENBR/C(?GRP 1���Cz  A��# �!��/�/�/�/�/ 6!
??A*ՀUr(A!~a+MSK  u%4}1a+N.!%[�~2�%��?��VISCAND_MAXs5�I�](�0FAI�L_IMGs0`����#}(�0IMRE/GNUMs7
�;BgSIZs3&����,CONTMOiUQ u4��PE���c�� �@�~�"FR:\�?� � MC{:\RC\LOG�F7B@� !�?�O��A�O_�z �MCV�O�CU�D1*VEX3[��`�qF�"ᖉ�`(ޣ�=��͍_�� Z�_�_�_�_�_�_�_ oo,o>oPoboto�o��;PO64_9C��B ��n6�eK L!IA�j�h�aV��l�f@�g�o� =�	�hSZV�n�����gWAI�o�4S?TAT �+�!@�O���z$����5J!2DWP  ?��P G)����a�;@'��2_JMPERR 1㖋�
  ��2345?678901|��� ����ď��ɏ��� �B�5�f�Y�k����<N0MLOW{~�@�0ζ@_TIYH�'��0MPHASE � %���3SoHIFTO21"x[
 <���?\�� ;�a���q���Я���� �ݯ��N�%�7��� [�m�������ɿ�ٿ �8��!�n�E�����*	VSFT�1�cV�0M�� S�5�q� � ��E�A�  B8������� p�����ª��B ��ME$�u4�q���a{~&%���M��x[�p�30��$xpTDINEND]H^8t�Or0U?�ׄ[J��S�ߏ���s5����Gy�	��,���������ߍ�RELE �s/q�XOjFt�?_ACTIV��~8<��
 A �;}�<���RD�`��C!YBOX ������v��p2���>�190.0m.��83����'254�����`�� �q��robot�ę� ?  pHa�upc���u���p��r���ZWABC�#�-,u�  �r�5X?Q cu�����/@�0//)/f/�Z;D�q���