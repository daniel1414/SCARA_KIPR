��   �A��*SYST�EM*��V7.7�077 2/6�/2013 A� ���$$CL�ASS  �S��(��D��D VIRTUAL%�7MNUFRAM�E AF�D� � 	� 88�?� ��}��y���� ��1=gQ s������	/��/?/��WNUM  ��>l�  �WTOOLa4� 
wN%M/��C� 3/�/�/1/	?3???? i?S?u?�?�?�?�?�? �?O�?O)O+O=O_O��OsO�O�Ok(�!{&
���&* 