��   D�A��*SYST�EM*��V7.7�077 2/6�/2013 A� 
  ����CELLSET_�T   w�$GI_STYS�EL_P �7T  7I�SO:iRibDiTRA�R��I_INI; ����bU9ART�aRSRPNS1TQ234U5678Q�
TROBQACKSNO�� )�7�E�S��a�o�z2� 3 4 5 6� 7 8awn&GINm'D�&��)% ��)4%��)P%��)fl%SN�{(OU���!7� OPTNA �73�73.:B<;}Ta6.:C<;CK;CaI_DECSNAp�3R�3�TRY1���4��4�PTH�CN�8D�D�INCYC@HG�KD~�TASKOK� {D�{D�7:�E�U: �Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T�8�T�@REQ�d��drG�:Mf�GJO?_HFAUL�Xd8�dvgALE� �g�c�g�cvgE� �H�dvgNDBR�H�dg�RGAB�Xtb�  �CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVIRTUAL�i{q'61ION � ��1��q�t+ UP0 �u��qStyl�e Select� 	  ��r�uR�eq. /Echuo���yAck����sIniti�at�p�r�s�tH@�O�a�p���	��V  �����������q����𱇪q��sOpti�on bit AJ��B����C��Decis�co�d;��zTryou�t mL��Pat�h segJ�nt�in.�II�yc�:��Task O�K!�Manual opt.r�pIAԖBޟԖC�� decsn ِ��Robot i?nterlo�"�>>� isol3���C��i/�"�z�ment��z�ِ����~_�status��	MH Faul�t:��ߧAler���%��p@r 1�z L��[�m�+��; LE_COMN�T ?�y�   ��䆳�Ŀֿ� ����0�B�T�g�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼�������������U������   ���ENAB  ���u�����x���ꐵMENU>���y��NAME ?=%��(%$*4��� D��p2�k�V���z��� ����������1 U@Rdv��� ����*< u`������ ��/;/&/_/J/f/ n/�/�/�/�/�/?�/ %??"?4?F?X?j?�? �?�?�?�?�?�?�=