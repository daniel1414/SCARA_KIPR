��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARA�M  b��ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
  ��APCOUPL�ED1 $[P�P_PROCES�0 � �1�V��UREQ1 �� $SOFT�; T_ID�TO�TAL_EQ� �$,NO/PS�_SPI_IND�E��$DX�S�CREEN_NA�ME �SIGNj��&�PK_FI� �	$THKY�P�ANE7  	�$DUMMY12*� �3�4���RG_STR1� � $TIT^�$I��1&@�$�$�$5&U6&7&8&9'0''�%!'�%�5'1?'1I'1S'1�]'2h"�SBN_�CFG1  8� $CNV_J�NT_* �DAT�A_CMNT�!?$FLAGSL*�CHECK��A�T_CELLSE�TUP  P�� HOME_IO�� %:3MAC{ROF2REPRO8^�DRUNCD��i2SMp5� UTO�BACKU0 �� �	DEVI�C#TIh�$5DFD�ST�0�B 3$INTER�VAL�DISP�_UNIT��0_�DO�6ERR�9FgR_Fa�IN�GRES�!Y0Qy_�3t4C_WA�4H�12H�W~0�$	Y �$DB� � CO5MqW�MOJWH�.
 \�VE��1$F �A��$O��D�B�CTM�P1_F�E2�G1Q_�3�B�2�X_�D�# d �$CARD_EX�IST�$FS?SB_TYPitA?HKBD_S�B�1�AGN G� �$SLOT_NUyMZIQPREV���� �1_EDI}T1 � h1�G=H0S?@f%�$EPY$O�Pc �0LEToE_OKRUS�oP_CRQ$�4x�VAZ0LACIw�Y1�R@Pk �1w@M{ENP$D�V��Q�P��A��nQLv*OUyR ,lA��0V1AB0~ O�L]eR"2CAM_�;1 x�f$ATTR�MP0�ANN�@�IMG?_HEIGHQ�c�WIDTH�VT�C�U�0F_ASwPECQ$M@gEXP;�@AX�f��CFT X O$GR� � S!1z�@B`NFLI�`<t
UIREs3��tGITCH~C�`N�.0S�d_L�`�CL�"�`EDkp;tL0J*DS�0>0�zra�!�hp;G0 � 
$WARNM'@�f�+P� �s�pNS=T� CORN��1�FLTR�uTRA�T@0T�p  $ACC�1
� ���ORI	`!S<{�RTq0_S�B�qHuGI1 [ �Tpu3I8�TYPVD+P*2 �`v@�� 1R*HD�cJ�* ���2��3��4���5��6��7��8���9��qO�$ <� #5x�s1�v`O_M�@�C �t 0Ev�NG��ABA� �c��@YQ������@������P�0����x�p�PyP�2� h����J�_R���BC�J��2�J	VP�CR��}@w��lu�tP_}0OF� �2  @� RO_�����aIT8C��N'OM_�0�1åq3�FCPT Ԑ#���@xP��J}E!X�G�0� .��p��
$TF`��C$7MD3��TO�3&@yU=0�� �)H�2�C1{�E͡� vE�uF�uF��0�CPo@�a� 	P�$@`PU�3�fc)"��)�AX 1�rDU6�$AI�3B�UFV��o@�! �|�pڶ�pPI�U�PZ�MY�Mf��̰i�FZ�SIMQS��/��A-�������kw Tp{zM���P�B�FACTqbGPEW6��Ҡؕ�v��MCc� �$}1JB�p;�}1DECGڙ�G��'��b� ě0CHN�S_EMP��$GO���+P_��q3�p2�@Pۤ��TC��{r ��q0�s��a�/�� �B0���!	���JR!0��_SEGFR��Iv *�aR�TjpN%S+�PVF�����ʹ Y�K��a1�)B��>�( 'j�Av �u�ct��aD�.0���p*�LQ��D�SIZC������T��O����>�aRSINF��� ��jq��C��C�����LW�����x�CRCLuFCCCkpy��� ��N}���bA��������d��DwIC��C ���r��+ P��z�2SEV2�zFH_�եFpNt/�>�,���H�1Q��!  ��@�Qx���� U�kp�2 ��a��s�+���A��S!x �"�4�4u2��tARt���`CW�$LG�p��B�1�Pr�P�t�a!A?@z�ϣ~0R���ME�`8�oC�3RAs3�AZ���4�pb�OS�FC�b�`��`FMp�� �0��ADIS+�aV%��b��z��pE$�pRp�cV�S0�P��a+QMP5�`IY8C��Me�pU���aUS" $=�TIT�1�S�SG1���#�8��DBPXW�O! T#��$S�K��2�P
0TmTKRLS$l�Q0TQ���P`P�D�q�1LAY_CAL�1�R^0�o f7PL)A�Q�D�'a�73a�7���AD�B!S%2?�PRj� 
*0���Sg& =�A$��S$ �*�L�9'�?H'�U�T(ODCS9)#ODENE��c*BO'Ӳ0RE�p�B+H �O�u�&$L�C'$@�3R��K2�LVO�s_D~!U�ROSbr�q�v�R����CRIG7GER�FPA�S��>6�ETURN�B�c�MR_}�TUbp\���@EWM$���cGN=`���BLA���TUܡ($P�')$P s�*hP3ab��C�TΣ@DO>����D�A���FGO_oAWAY�BMO"��a�!�DCS�_P,<aIS t�� �� �s�S#�Q���Rw�cV��Q�w2�VW��'dNTV(��RV;����~��mgŃ��Jt��<@���SAFEڥ�f_S}V�bEXCLUT�:�� ONL���cqYfЀ�y�OTEu�HI_V} ��PP�LY_�q7�VRF�Y_b3���Rj L�_G -h@0��_y��1� ���QSG�  .�rŐ1PNQ�5�� _q���;P��V�by|rsvANNUNX<@�$�tIDX�UR�c[P� �y�qi �zZ�vT)1EF�PI<B/��$F�r�$А�OTQP�A $DUMMY��&����&���*0t�U0 7`  �HE�\����^r�cYRr SUFFI���Pa0���P)�5#�6#��DwMSW�U1 8���KEYI��4�TM`�A��ځ3QՆINݱ�v�
)1j P2 D���HOST�0! ��������������EM&����*0S�BL� UL��3 AZ���D�*0T�@~S4 � $���USAMPa༥.������V I�@��$SUB����;@�c����3��SAV �����������`��vP$�@EC!	0YwN_B35 0��DI�t�PO\�M��#�$E�R_IB�� �ENC2_S��T6X��2������� �cG���0 S7�2��1��A����8  ��Ǜ��@�PK�Dk!uq��AV�ERҁ�����DSP�ܢPC?���2�6�\�����VALU��HE �M_�I�P(�ܣOPP� �5�TH��ͫ��SH` 4�.�FB�6d���~�� �BSC?q����ET�9ȂF?ULL_DU���q�KP�ԝ�����OT��"T�PNOAUT5OS:�$YĪ�Z� ���X�C(02h�CE26p�V��L� ;H *h�L� �����$P��wc�ě1�Ʃ1���C��Ƨ��Ʋ���7*��8��9��0����U1��1��1	�1�U1#�10�1=�1Jڥ2X�2����2��2�	�2�2#�20�2�=�2J�3X�3��3T����3	�3�3#�U30�3=�3J�4X��[���SE�2< A<8�Z����I��0e�$�}�"qFE5P?P�T= ,f��a?3 �P�?i��Je�i�E�Pq�N��`T>F�$T�P$!$VARI�����UP21p? 7���TD��s���p�������q��BAC2@ T����$�uP�*��Þ0� IF�Iw�0�P� � )P�B"	N�0P�TAt ;u�"�"pu STvt: �btP�@�l�6	sC2	>0���S���/b�F��FORCE�UPsr��FLUS
�pHfNn����b/D_CM�PEv*IN_t�e`�REM� F�a�a��0�Te�KdN~�eEFF�j�PsINJa�OVM��OVA�TROV���DT	��DTMX,A��P*���0M(xR#�0�CL�*_��u*�Pr�{_�XЉ_T�+X�J�PASaD% ��(�װ�1`�&_A@RQ~�LIMIT_�d4�� M��CL�t�ˑRIVW�*2E�AR�IOxPC��P���B�R�CM�QP*�b !GC3LF�#�1DY�8} l�q�35T�%DG�h��0�5+N�SSt0��B P��1�A�E�`_�1�8�11���E�C�13 K5 F��GRA��gC��4k�`W�ON��"EBUGwctBx#p�C ��_E D ����`���TER�M�EE�E  ��ORIS�@F�F �SM_�`���@�G�EԠ�TA�IHܙE�P�UP��Ig� -�Q��D|`|�C|PE$SEG#Zv�0EL�eUSE�PNFIzLRT�kAx,��DTF$UF�`O�$\��a�P/���Wi@T��t �cwNSTTPAT��<h��RPTHJKa-�E
�65MR<p&�WUw��&�Q�LQR<`�Y�qS�HF�pYT�Q�X_SGHOR�*��F �@�$�GM`H�u OV�Rq��q6`I`4Uz� �aAYLO���"J�Iu2b��Q��o���ERV���a� 6j �WnP�R~�E �e���E Rb1Pp�ASY1M|�p�MQWJ`W�� E���Qy�b0�U�7tnPI��Uw�/�eP�o��`o�fgORnPM|�S�GRSMTf�Jg�GR��aC�qP�A|P��p=��K ׸ FTO�CFQ�P9`N $OP@/��#��N e�!O�ڐRE
��RdS�QO����Re�R�UN�%�a#�e$PWR0IM@��bR_ ���=�mR� LVBH�_�ADDR$�H_LENG�Rǁ���T�uR� SO�M H�S���~�����Ì�	�SE!u���S�:�MN�1N���p��F¹�OL���8�3�3�=��ACROc�z�P$��[�p�a;�  �OUP����r_�I���q�q1 �ѭʓ��ԙX!՘Y1 ՘t!՘	�ԙлE"IO���DϗA�ߕ<9�gO $���p�)_OFFb�;�P�RM_Ò�qT�TP_[�HjP (��OBJ�2��#[$$�LE�S��>�Q � ����AB_�!T���S��p;x LV��KR�32@�HITCOU�BGE�LOہ 磴!��@��"�G#�3SS��HWD�SQ�jR�lpINC�PU��VISIO �����Ğ�
������~	� �IOLN�S� 0C$�SL�r@PUTM_�$@��PV0x�ɱ)F_AS�2T $L  �� D=a0U�@9`dQٵ��䳊`HY#�]�6Ù���UO�3U `"�{�$�5"M�5 Tƥ�R�P;@��ǿ�hT��µ��UJe�V]���NEfgJO9G{W��DIS��1K��� �3W XХQqVv��P;�CTR�S�:�FLAGBB�LG�tX �� ���~aCLG_SIZ�����d �����FD��I�اؓ�׏ث@ �֎����	�d 	���	��	�@	�% SC�H_��R���aBg�NTє�Y��!E�2��p�J U}�}��p�L��|�DAU��E�A�����t���GH��rf�OGBOO>Zh A<�f0�IT2���@8�REC�SCRB�=��D:�����MARG �<18��0��a�%�Sȣ$�W?�%����0�JGM��MNC�Hz%�FNKEY���K��PRG��UqF��g`��FWD���HL	STP��V`��mP������RS;	Hp��-�Cid6r0�.0s��	U|���r� Xb��P�E���G��`CPO�
.�M��FOCU�RGE]X,�TUI��I��p�K|�V��V�� ��A`B���p�A`�9Nu��SANA%�FRޚ�VAILy�CL�P1uDCS_HIyD�
��O�X1��S� ��S�V�I�GN��~�ӽ�\�T|���_BUFF�1�[5�o`T�$ ��� ����B�`R"�
�1\5�o`ܰ��c���pOS1�%2�%3�!����0] � ܩ�qEU������IDX�tP�bD�O�� ��Q6ST|�R��YV�@1 \$EO6CO;�{�^6�q6�%��0^ L ��K�[@`�9`(��S����:�����x��_ _ �pp�Ð���� C�@Cp�` ��� CLDP|�uTRQLI��Ft
�4I"DFLGV�"@1VCb�D)�VGr�LDVE@DVEORG
�qiB _�g�H
��d�D�ta �0�@Dr1DVE�S�pT4@I��@T>VRCLMC%T�O0�O7Y�� MI��tgb dy��!RQI�=0�DSTB�0c �VO�XAXr� �X�\EXCE�S6�t�vRM_��qc6��Rt��vR<��p5d��V_A�Z���(k�_�X@K�te q\����/�$MBs��LI���cREQU�IR�b��l���hD�EBU��sQL�0M,�f�r��`����%R�sQND���p�pg0w�n�?�sDC��IN����p�,x' �NV���K����bP�ST� h��L�OC�&RI���%E�X�vÀ�!�QsQOwDAQ,�i X��3ON���MF\��� �v9�2%��5�uk�0��� FX�PIGG>�� j �M��2�!���3��4R �%?3;�|�K�|�Z�G`�E�DATA{'��E��U��b"���NZ"k t $MD��I��)Ɔ ф��ф�H�p�`Ѕ�X�҃ANSWe�ф�!'х�D[�)�r��P��l[ �PCU��V��X@�uRR2��m �D���a���Rd$C'ALI�P"�G�w��2��RIN��z�<Nu�NTEڰ�"nI�`��°r��ڰ_N���oÕޒi�oT۔bpn�DIVmVDH�Ptݐ��q� $V���+s1$��$Z �"��� �"f�_�e��rH �$BE�LT>��1ACCE�L!������IR!C��P��t�T31h�O$PS�P'BL� M�ʤ<C���������PATH�����"�3ТZ��Q_�!U��2�8�R� C堌�_{MGP�$DDU�<��/�$FWh���`��q�����f�DE���PPABNاROTSPEEH��!��4@J��!��P��� ?$USE_���P��O�SY��g�Q- B�YNyPAO���OFF��MOUfR�NG�O�OL�L�INC.��q��u��Rn�PP�RENCS������Rȡ���TŠIN'2IТ���`R��VES�{���23_�UPI���LOWL�!� �4@���D�� �R{`���0��5bC�ΐ��MOS4 LdM�O���PWPERC7H   �OV�� b��!m�@1�^T@1�s@��hP�`�� V5�'`ѡ��L���Ig�Ԇ��UP�Ӛ���T�RKv�#2AYLOAA��$a1�Т@�5�8�p40��RTI(a|�40MO����R$b�@N��T��w�L���"�f�DUM2,�S_�BCKLSH_C Т��B�A�u�'�Y��������6�x�aQCLA�Lz ���Ar�`�C�HK4@+5SH�RT�YS��}%�A��_�:36�_UM(`n�C�{�c�SCL��ʰLMT_J1_LS�"�P������E������������SPC`��;���	��PCs�B��H�0�`Y�q�C3P��2XTc�g�CN_"��N��i��SH ���V	�*3�Ň�=Тd�AC� y�SH:3 ��g��ƝA���s�4�0ѡ��c�PAx�l�_Pw�[�_5@��8�`V�4AH�ZK�JGG"�M��OG[��TO7RQU��ON.�Q����wbLҠᝰ�_W��1�_A��G��M���I�I�IM�F��p�JPQ2(�A_�VEC��0�T�RS"1Y.p�Pm/�R`%JRKY,��"�&PDBL_S�Mh�RM)p_DLG�RGRV��$G��$M��!H_ �#��:COS;`�8LN� ;;\%B4G�=9M�@=9!y:g<-!�%Z60�L־!MYD1�8$2T�H*=�9THET0�NK23M�BA��E0CBFCBA�C �Q�R,B$:AG�:AF�SBG�XBEGTSaʱC��qW4&��Dg3�Gv3$DU H�Ih�Aw�x��R�F��r�QQ���v$NEd��IF0Y�`R�E��$%��1A�5#U,W
581LPH(eR��RS\%tSg5tSv5R�6P�S�Z�6%�VEXV:XT7�]\VlZVy[V�[UV�[V�[V�[V�YHEX^Vdb\]�{hy[UH�[H�[H�[H�[UH�YO6\OEXO�i�[^OlZOy[O�[O��[O�[O�[O�6F�R'A�yg5�t8WSP�BALANCE_l�1�sLEo@H_�5SP��X6�rg6�rv6PFULC�x��w��v5Ț1n}�UT�O_C�nT1T2G���2N*�z���g����k���@ע����T���O����INSsEGz�%�REV���%���DIF��1�o҇�1p�pOB0ȁ��#��MI��5�~�$LCHWAR��悢AB*y�$MECH0A�0>�D�Y�AX>�P��]�W(�<�q 
^������7ROBV�CR�Ҡ�zR��MSK_�p�j�s P R�_���R��H�Ҕ��1 ���ԲҐ����Ґ&��IN���MTC�OM_CD n�t � P�ڀ��$ONORE��9����(�u 8�GRl�I�SD�@ABJ��$XYZ_DAx9Q���DEBU��XM��U�v �p$�wCOD�� ���o�J�j�$BU_FINDX԰��MORœw $1�U��-��v�F�����Д��Gܢx �� $SIMU�LX�����$���O�BJE�p$�ADJ�USB�5�AY_I�o��Dc����G�_[FIJ�=�T� ���������������Հ�P��D�FRI4��׵T��RO����E�����OPW�O� ɐy0��S�YSBU�PΠ$SCOP���#�'�U&˞ՀPRUN�M�P�A�DL�H�!���_�OU�!A���r��$��IMAG��4ϐ�@P��IM�����IN� u£�RGO�VRḎ>°Ѐ�P0����԰�@L_:�����m� RB� �@2M��EDՠJ� ��NpM.�������SL�pɐz x $OVSL��wSDI��DEXq@k�i�=!{��Ѕ�V���N�Ѵ{��Њӟ�Ěط�M�!РF�_SsET�ɐ{ @����g���RI&���
��_4A��	����ׁ|@��  | Hϑ�I�J�ATUS��$TRC�@ǰˢD�BTMM�7�Ij����4��#�,�ɐ} �DϐE~�k�A�`E�ۂBᏱ
��B�EXEH�Z�ќ��{���1~��АG�UP���s$����XNNm��=!p�L!p� �PGn&��!UB6��g��6�
�JMPW�AI� P��N�LO��j�F��#�$R�CVFAIL_C�j�Q�R��Q�Z�M�� 𣕠���0R_P=L
�DBTBm��j�BWD��A�UM���IGe���m�� GTNL� ����R���.�Ep�һ�!��DEFSPy� G� Lϐd�7 _: H�HUNI��r�F b��R��^�� _L��5P@����P�ȑ����F����Ѐ��p:��N�pKET�}��� P��ȑ� h~W�ARSIZE���l���S@�OR~
�FORMAT3����COJ����EM2V�lUX�����PLI��ȑ� � $#�P_S�WI�i�%��AX�����AL_ ���E A��B�,@C���Dj�$E����uC_��	� � � ���q�J3�@����TIA�4�5�6��MOM�������#�Be�AD�&�&6�PU;@NR�J%��J%�DŔ�� A$PI�F�ޑ ��$�%�#�%�#�%=D��&�+QD�DpсF��U���g�SPEED�`Gd*4f�716 7f���16g3@8��8O9��f�SAM�p�p�417�3f�MOV�� �D�1ƀ�E�4�E�17 	1��42��������5n��Hm��3IN 2Ln�39HUK0Df�;J�{HRD{K�KGAMM��v�A�$GETH��ȠL�D� �
b�OLIBR��I��$HI��_��P��bVE�XA^:P+VLW]XVO\:Y|V+V�V����� ?$PDCK�U�"L�_�0�� �.B� m!E�W��T&�Yr� �$I�R�S�D��&����(�L�E�ޑ�Oh�)`�qE�ɐ�P��?UR_SCR��a�^��S_SAVEc_D�īe��NO�C����`�D��& �i��)�iapz{p ���&Ex@�q��0�B ���5G�2�+8!�;6���g8�w�ucs�1��:EM{%� ���� !G����c�w���`ζB�qW�`��$��0��N ��R�qM��H�C�LG�GM�aǒ� ?� $PYr�g$Ww�+�NGt� �w��u��u��u� �������@[L�n%X� O�mZ��GQ�Ŕ� pW�#�c�&�o�o#5�:�_)�� |Wи �`��������`�ޗɖ�EQ��EB��J�b�Ϡ���P���PM��QU�0 �� 8� QCO�Uas�QTH��H{OL��QHYS3ES�1[�UEG��b�� OM�  �P�4�U�UNI�J�� �O��)�� �P�������a��R�OG�j��2��O�𤥥c�󠉠INFO(�� ��ث��
��1OI�� =(`SLEQ"6D� 5D�ܦ����DS𿠉���VPO�P�0#3�QEMPNU����A�UT�a��COPY��1�಼��`M��NH������CT�� �_RGADJ(���X#�_$� '��
'�W%�P%�]`'�:3l�;�EX��YC��I1@OՐ(���n��_NA�1!S����i����M� � ��p�PORp��Ì&��SRV���)����DIT_ p��� ��
��
�w�
�5�6�7�8���1S�b�����M�C_Fe��pL�a�a�;�Rq���/��җ#�0��k��� ,`FL����`SYN{���Mp�C���PWR���������DELA �6Y֨ADR��QSwKIP{%� ���Z��OŀNT�1�p*�P_����I�`߂ ̐`��#`�3`��n� kn�;�m�H�m�U�m��b�m�98a�J2R�.0��� 4� EX�@TQ����q����������jRD�Cx�� ���X��RF�E@AY�_�X�~�DRGEAR_�@sIO�t=bFLG����EPC��U�M_���J2TH�2N�# � 1��UA�G�@T�P I�"���M��-�I����4,��REF�11�(�� l!�ENsAB� ��TPE2` {� 8Wܠ�M�q �CL��R�w��2'�-?Qcu��3'����P���4'�'@9K]o��5'��������6'�!/3/E/W/i/{/�7'��/�/�/P�/�/�/�8'�?�-???Q?c?u?�SM+SK(����� �E�axaREMO[TE���
��`0/B`��q-CIO�UQE)I�0�R� W\`��� /���-�����ҿ���ՈB$DS?B_SIGN'a�qĘ���C��pS2�323E���$�DE?VICEUSKC�r>�rPARIT!�A_OPBIT�q��OWCONTR����q�0�rCUPM~�sUXTASK�S�Nq��P�DTATU��ppBS3`����u�e�_�pC��$�FREEFROMqS������GETA`.��UPD��AEbfS�PTP���� !>�8$USA����x�9h�{�ERIO��L�`ՐRY�U�B_�`��P�QQfWRK��?�<Dh�3fh��6F�RIEND�qg��$UF�U�p`TO�OLwfMYd�$�LENGTH_VTߤFIR��cM��SE�@�iUFINttrаARGIa�F�AITIi�gX�F�i�fG2�WG1`�� �Sr$wPR��sau�O_�@�P��xQ�RE���SU�ءT�C�N�=qyv �G(��]R���u��Q�A ��hzhZUz�ZU�t����{P�T�X T�P��L��TcH���hh�U�T�SG��W$X�)��r>�D����.��C�z�N�b��=$�v 2�!�-a�' 3i1?h.`21k2
��31k3?j���@i�����6{��s{��r$)V��bV�eV���vYr���O�[V{�@���hv3Ru�^pib��P5S��E�$���c��5$A8й�P!R)��u,�S���@���V�¯ 0�p�v���P�N�����!��P>p ��
�US^zA� �\�R���GA_�Š��Ny@A)XQ��Ag`L�ag�^p�THIC'a��8-����QTFE���>m�IF_CH'cp�aI_����6D�G1՘�٤*��h��`��_�JF�PRW�I���RVATF�� ��\�'�f`��)�DO��e)�COUW�C�A�XI�D�OFFS=EZ�TRIG�sz��,�)�#g���z�Hx����g�IGMA�P��a\���ȸORG�_UNEV#@Ͳ ��SD���d ӎ$����GR3OU[A�TOa�Q��DSP#�JOG�V�S8�_PV�3RO����U�mpEVKEPF��IR?�_�=pM �&��AP���E�������SYSv��B��;PG��BRKYr����b�\���������k�ADVQ�y�BS�OC�C@N�DU�MMY14��`S}V�DE_OP1S�SFSPD_OVR���C~�N�QÓOR\׶0N�P]�Fء�]�<�OV?�SF��a����F���Ac��As�؁a�BLCHD}L�RECOVM��P<�W�`M<��?�#RO1S�K�_a�_�� @���`VER�t�$OFS�`CV�@_bWDv� �rѰ��R��9�TR%Q|A�E_FDO�ƟMB_CM[A��B/�BLl�_¦�l�甁V�qDb�P����G���AM�Ú�yP��'��_M��>R��HC4�8$CA2���Ȱ>��8$HBK�Q��N�IO1e]�iAA�PPAQ�}�b���u���iB4�DVC_DB�c�񓡦B����A"��1��'���3��-�/ATIO�@��FP�M�UDc1�HFCAB H�0bFs�p�p��Ea�<�_BP��SUBCPUk�I�S%��@�� ��P�s�,���B��?$HW_C!���i��x�A'q\�l$�UNIT��l�A�T}����I�CYC=L��NECA#���FLTR_2_F�IҤ�H)�FEaLPxU˲���_SCTosF_�F��
v�
�FS�A���CHA�Ja^���3R�RS�D1�B ё�l�i@_T��PRO ~�)PKEM�0_���8��3� �<�*%D�I�P��RAILAiC��rM��LO��c+�i���-��-V'�PR��S{q�0ҕ!C���@	&�FUsNC�³�RIN�p`Z�+`? �$(QRA� mr 9��#��G��#gWAR�:�BLuq��'4A;88D�A���!I835LD@�PA�A�q3h��!��q3TI���5�β�pgRIA�Q�BAF� P�A���1��5��T����EMJ�I1Q��D�F_�`�ӨQ��LM�t�FA�`HRDY4d�P�`RSoq+`|Q0EMULSE�`x���E� ���I�����$]a-$�Q$�Q�,���� x��EaG�@�AРAAR�2)�09mb�E50��wAXE&�ROB#��W�ac�_�M�SY����Ae�VSWWR�ذ�M12�� STR�"Ņ�d�h�E� !	CUq#��lqBhP3�oV��)��OT�Pv� 	$�ARYg�ЦR_!�`	T�FI���j�$LINK(�1w��Q�_eS3��CU��RXYZ@Q��[��	co��Q�RJ�X�PB!��"Kd0�
 � LcFIeg`3�D�9Ԫ$<�_JN�p"�e��SA�OP_~T2�[53�NqTB�aNB2�bC9��DUQ�BV=6r%TURNb����u�Q�!h�?�gFL�)���B�@+pekZ7�3�I� 1�nPKH�M��BV8r%����c�ORQ&�!�# mX�C�����갦��up��.�<��tOVE�q��Mj�tC�zC��B�W�Fq�� � ��� j�0���qw�P� ���	��q���zC��L5��!ERM��!	v"!E8P���#؄A���id�%"�WP1MP1AX�bP1��&!�Q2� 2!>�\A>���=��`=� p=�ep=��p=��@=� JQ=�@:�@J�@Z� @j�@z�@��@���@��@��ב˙DEBU�$�!�1($�{�P��R�g� � AB�P'N�[��sVְ� 
����Ϥ��Ϥ aڧ$aڧ�aڧqڧ eqڧ�qڧ�A�4�`�2\�RLcLABbb�u� ���1s  ��ER�9P �� $8`� A�!��POB�FЉ�P��ލ�_MRA��� �d O0T<�\�EcRR:�2�0TY��aIA�Vb`,���TOQ+�i�L�@,�7R����� C�A � p�T�P��< _V1ْ.�V�2#cą2\�2k�ȱ��op�8ˠȱu�$W��j6�V�A���$�@"�0,���6�Q�	�@�HELL_CFG��A� 5e Bo_BAS��SR��\p�� �CS�T�1�1��%�22�U32�42�52�62�e72�82��RO ��8��P,`NLzA�cAqB��H �ACK�� >�i���`�`G@���7_PUr�CO�@��OU��P0�W!���3�7LTPX�_KcAR���RE���&@P W1�QUE�� �p9CCST?OPI_AL������PU#�Д���PSE�M���M���T�Y��SO��W�DI�����}�L�1_T}M�MANRQ���PEZV�$KEYSWITCHU#�8��CHE9BE�AT!�E�@LE(�$f�U4�F��5�|K��O_HOM�0�O�#REF�pPR��!)�AUP��C��Op�0ECOư_1`_IOCM�d����S����g�@� �D�Q� U۲{�M�w2Q��p�cFORC��3 �@��OM>�@ � @���3*�U[SP�@1��$��@3�4�1��N�PX_AS�¼ �0�ADD' h��$SIZ�$VsAR2�D@TIP��)�� Ah�аJ� � �� �BS��AyC��%FRIFa���Se�w	��NFp�@Џ@� x�SI�TEFsj"es�SGL}T�R7p&�A���#P~STM�TJ�P�@;VBW<�pSHOW�R���SV
@�D��; �ԱA005pЁ  "� '� '� '� �'5)6)7)8
)9)A)�@'v  'V�	&r`'F(JP �()�P�(,)#`�(F)@p�(`)�p�(z)1�)U1�)1�)1�)1�)U1�)2)2)2)U2,)29)2F)2S)U2`)2m)2z)2�)U2�)2�)2�)2�)U2�)3)3)3)U3,)39)3F)3S)U3`)3m)3z)3�)U3�)3�)3�)3�)U3�)4uI4)4)U4,)49)4F)4S)U4`)4m)4z)4�)U4�)4�)4�)4�)U4�)5uI5)5)U5,)59)5F)5S)U5`)5m)5z)5�)U5�)5�)5�)5�)U5�)6uI6)6)U6,)69)6F)6S)U6`)6m)6z)6�)U6�)6�)6�)6�)U6�)7uI7)7)U7,)79)7F)7S)U7`)7m)7z)7�)U7�)7�)7�)7�)�7�$%��VPd�U�PD��  ����)и�YSLO>��� � ��0�Q��TA�����ALU������CUT��F��ID�_L��HI�I~V$FILE_��?�+�$��SA���� hҰk�E_BLCKh�x����D_CPU��� ���� �B�T���q�	�Rw �G�
PWl��� �LA1Sp������RUNu� �����8�u�?����?�� �T?�AC�C��X -$f�LEN��s����f�����I�J�LO�W_AXIh�F1f�,�2��M��	�G��_��I��Y�8�թT#ORn�f��D��ܣ\LACE��Y�f�8ٳY��_MA� ��83�	�3�TCV:�[�	�T�\�{�q�|�������	���J����MDĴ�J9�����
	�r�2�Ц�����l��ΠJK�VK��h#���#�3�J08Ķ'�JJ/�JJ7�A�AL'�]�/�]�W�42X�5��{�N1����(M�I�ڤLӠ_���Q b���� `u�GROU����}Bd NFLIC���REQUIRE��EBU��b�Ŷ��2�c�	�a�� ��� \APKPR�C �ܠ
a�;EN\�CLO��lهS_M`������
�a��� �F M�C6�{�����_MGV��C�l��؎�5����BRK��NOL������R�_LI��������J��P _��/��7��{��D���6L�O�8����>��� �ҍ�z��燡��PATH�������ᒨh��� $��ͰCN���CA �]���INFe�UC٠��%�C��UM.�Y��4���Ez�P���P�7�P�AYLOA�J2=L��R_ANE���L���������R_F2LSHRC��LO��$���2���>2�ACRL_�"�� �����H�b��$H��CFLEX�_�`�Je�� :r���	�t���`��	�������F1� ��ïկ�����E'�9�K�]�o��� �������$��гĀ#(ؿ�����TR'�X ˲�`H ��%�&�8�J�\�`� i�W�{ńϖϨϺə�}J��� � ��0����ʁ��AT�6ðELt �5صJ����JE��C�TR�TN"F��6	�HAND_V�B�_����� $f F2�֋���SWF������O $$M���R�Ӏ�H�ѕL��E:�FA@�������I��A��݀��A��A	��@��T����D��D	�P��G	�qYST��yQ��yQN�DY �Z��� �D�E��)��������@���H$� � �PT� ]�f�o�x����}3>�� {@`��n�xvf��o�ASYM������Ͱ����_SH��#�=�'��dLHG�Y�k�}���J���G��gs]y��_�VI/C�x�ӵpV_UNI���t�#��J��re�r���t�� �t�ð	G�(:�j��#PXI��TA�H��N���EB��EN/@��DI	�W#O���ᙀ�ç� � �BI�aA K����吂��U��0�`��n�� � ]AME\?0�g��aT��PTpi0��5�����K�,p:�U��I�TKp�� $�DUMMY1�!o$PS_RF� �  ����͑LA���YPV#��=�$GLB_T~@��ŕ�5���`�CAӁ� �XI�	נ�STȱ��SBR��M21�_Vɲ8$SV_�ER��O��#�C)Lߐ�AuO炔���0O� � D� ĐOB���3LO�f�S�y�ÐS�p��1SYSS�ADR��1��5�TCH�@ �� ,f L���W7_NA
�����y5SR>��l }J�J���F� �B���G���I���ID� ��D���D���V�p�KY V���bu���ݻ�������);Mt��XS�CREi�W��E@f�ST��F�}��La�Ǥ��0_�0AV�� TI�&��� �1%������1��ŵ��O�PIS�1أ����UEЄ� ��񪠞�SG��1R�SM_����UNE�XCEP��ј�S_ߑ��7��&�9�T���COU\ғ�o 1֤�UE���؂6�y�PROG�M@FL�1$C�U&�PO�>��I�_�H�� � �8E��_HE_�������RY ?��0���������O�US � @���D�$BUTT�/�R����COLU�M0��s�SERV<�3��PANE�0V�u��TpGEUA�|�F��ʡ)$HE�LP��bETER5�)��E���Oq��30 ��;0��M`��U`��]`���IN��-�TpN(p��0�131�o �i�LN��'� �0���_�����$H_�0TEX��3j�^�~$REL�V"D��~Ӑ�b���Ms�?,��p��4�򪑥#��USR�VIEWV�� <����U"�]@NFyI�0��FOCUA�n��PRI�`m���h� TRIP���m�UN��Є� ��`/��WARN|����SRTOL䥥�&�Rs�O�cO;RNsRAUW�v9T�	���VI�υ�� $��P�ATH���CAC�HV#LOG��LIM�r�S��BR'�HOSTǢ!����R|�OBOT�ƣ#IM� ��S ���0r��������VCPU_AVA�IL���EX�!�aN��} ~�Ma�UaL�]a ����{0�$BACKLA�S� �!�$"W�� � ��CT%s�@$�TOOLǤ$�_wJMP�� ���$SS�v4���VSHIF`у�PB���ǤЇ�R�k(�OSUR�3W�RADI�$��_���%�м1�ぺ���$LU�q$OUTPUT_BM��IM���b� }p����#TIL�'SCO�"�#C���$N�&N �'N6N7N#8�B��u%=,�2��0S �`Є�<��D�JUrU��P�WA�IT���<��:%�0NE~��YBO�W� �� �$������SB"IT;PEo�NEC/,B@@D(D�PJǐp�Rv @hE(�#=@�0�B�E/�M�KT���"y�� �An�!�OP�
MA]S��_DOآ�qT��D]����C��>RDELAY��SJO�"X֡�c'T�3���`� ��,l�y�Y_Ry�wR�#Ƣ�A�? G��ZwABC�� ��R��
Ȁ�$$�C�X�����Q���� �PV�IRT�_�PAB�S�!��1 �U�� < �Q(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�K�|`�AXLMTZvK��c  �]��INf�x�\�PREȏNk�����LA�RMRECOV ��Y�����@F {�UP   dK��"�4�F��T���w����������, 
#o�W�NG�u k	 A�   �,�`PP7LICu�?�U����Han�dlingToo�l m� 
V7.70P/36+�v�
��_SWr���F0���� 4�3�ˊ�yϋ�7D�A7�철
f���rm�None�����Oհ�P��T���<�_�+�V��R�v�7�U�TO�RX l���n�HGAPON�Pe� azn�U' D 1�� �и�����T��n�� Q 1� � �����P����	�7�H嵡]��R��R �a�,��H��B�HTTHKYV��R�+�=� O������3����!� ?�E�W�i�{������� ����/��;A Sew����� +�7=Oa s�����'/� //3/9/K/]/o/�/ �/�/�/�/#?�/�/? /?5?G?Y?k?}?�?�? �?�?O�?�?O+O1O COUOgOyO�O�O�O�O _�O�O	_'_-_?_Q_ c_u_�_�_�_�_o�_ �_o#o)o;oMo_oqo �o�o�o�o�o�o %7I[m� �������!��[���TO�C�U�DO_CLEAN��|5Ի�NM  	�Կ��+�=�O����_DSPDRYRL��HIa��@�� ��ϟ����)�;��M�_�q�������MA�X@���[����׳�Xࢄ���҂�7�PLU�GG�У���S�PRUCt�B�����Ğ��O�}�5�SEGF{�KY�k�v�� ����Ͽ���=�p�LAP����o�Y�k� }Ϗϡϳ������������1�v�TOTA�Lզ��v�USENU���� ���ߎ����RG_STRI�NG 1s�
��Ml�S3��
��_ITEM1��  n3������ "�4�F�X�j�|��� ������������0��B�I/O S�IGNAL���Tryout M�ode��Inp���Simulat{ed��Out��OVERR��� = 100��In cycl�����Prog A�bor����~�S�tatus��	H�eartbeat���MH FauylAler%	 U�CUgy���8��� ���� �����6HZl~ �������/� /2/D/V/h/z/�WORy��۲!&�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�?8OO0NPO�� V@�+?OyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_QBDEVYN�PmO�_!o 3oEoWoio{o�o�o�o �o�o�o�o/A�SewPALT �q�/x���� � �2�D�V�h�z��� ����ԏ���
��GRI����B��� j�|�������ğ֟� ����0�B�T�f�x� ������0�j�R� Z���� �2�D�V�h� z�������¿Կ����
��.�@�R�ԯPREG�~����dϲ��� ��������0�B�T� f�xߊߜ߮����������X��$ARG_�� D ?	����9�� � 	$X�	+[M�]M��X�n��,�SBN_CON?FIG 9�������CII_SAVE  X�����,�TCEL�LSETUP �9�%  OME�_IOX�X�%M�OV_H����R�EP�S�&�UTOoBACK�����FRA:\�x� Z�x���'�`��xǣ�l�INUI�px���l�?MESSAG�������A���ODE_D����#O�P2l�oPAUSVA!�9�? ((O<� ������� (^L�p���ej@TSK  �u����o�UPD�T) ��d ?W�SM_CF��8����%�+!GRP [2
5+ L�B���A�#�XSCRDv/!15+ �������/�/�/?? (?�����/p?�?�?�? �?�?5?�?Y?O$O6O�HOZOlO�?O(�r�G�ROUN S�CU�P_NA�8�	�r��F_ED��1�5+
 �%-BCKEDT-�O00�%_I_�� ���Q-r�_x�o�o�x���U2r_/��_�_�R�o�iU�_&o�_�_ED3o�_�o�_�n_o�o9oKoED4 �oro'�onn�o�oED5^�:�n����ED6 ��o��nK���%�7�ED7��^�����n�Z�ɏۏED8J�*_��N_m����m��ED9�[��ʟm7����#�CR_����7�ٯD��ū�@�@NO_D�EL�O�BGE_U�NUSE�O�DLA�L_OUT ���R�AWD_AB�OR�𦾦AݰIT_R_RTN����ONONSi �����CAM_PAR�AM 19�#
� 8
SONY� XC-56 2�34567890�H ��@����?��( С�Z���yŀ��\�HR5o��������R57����Aff��\�L�^�Z��ߔ� o߸��ߥ��� ���$��6��Z�l�a�CE__RIA_I(%5;�F�!{�x�; ��_LIS$��c%����@<��F�@�GP 1Ż���OK�]�o��.�C*  ����CU1��9��@��G��Z�CP C]��d��l��s��R������U[��m��v����}����� C���ő& ��G��;�HEנONFI���@�G_PRI 1Ż��T�������� �CHK�PAUS� 1I� ,�BTf x������� //,/>/P/b/t/�/O�����8�!�_MOR��� }��@2C3����<���" 	 ���/ ;�/.??R?\5�"�"���-=ֱ?99���3�@K�4��<P������a�A-8��?OO�J
�? KO�'ưS��"��:O��i`��PDB� ��-+�)
mc:c?pmidbg�Od�~�C:�  �P�P���Ep�O-_�C�P�7@�7@�V��@�Oq_<Z�.���.��S[_�_=Y�",�F,���UYg�_oV�\�װ�S[f�_�KoAMo�JDEF 3ch�)�B:`buf.txtqo��Mro�0����'�	z�A��1=L���j+MC�#�-,���(>ss�$�-�r���Cz  BHF3C�s7 C���C��M�F��iDP�E�~�WJ�I0D�tE�q�aEpIJ$��3HHƷ���{G�G���GG���N�[5K~w)L�{�XWI>��{,�iO�fu7��4�)�,�,�.װ�,�b,��@�u�K�x6�ʈq�* �* e�D��n��pEWLI0EX��EQ�EJ�P F�E�F�� G��}F�^F E�� F�B� H,- Ge��H3Y�WI�?��p�33 ��%WDn6��"��#5Y��\2��A�1WD~q<#�
 �O�+�)�Zj�bRSMO�FS���n6��iT}1� DE  �?fDR 
�,�;�&��  @�:��nTEKST�bo�8�R���!�/3�nvC+�A�WJq� [��rq��C�pB1 w�Cy�@�T�6��T�FP?ROG %ź��ů��I���𦶠喤�KEY_TBL � �6Q�!� �	
��� !"�#$%&'()*+,-./01g��:;<=>?@A�BC�`GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~�������������������������������������������������������������������������������͓���������������������������������耇�����������������������LCK�X	����STAT*��_?AUTO_D�����G_�INDT_'ENBK��"R��i��[�T2��\STO�P���"TRL��L�ETE����_S�CREEN ~"�kcsc���U��MMENU �1""�  <����|�WE[߅ߺ� V��߽�������,�� �b�9�K�q���� ����������%�^� 5�G���k�}������� ������H1~ Ug������ �2	AzQc �������./ //d/;/M/�/q/�/ �/�/�/�/?�/?N? %?7?]?�?m??�?�? �?O�?�?OJO!O3O��OWi;�_MANU�AL�Ϟ�DBCOƅ�RI�P�4�DB'NUM�`�<q*��
�APXWORK 1#"�ޟ+_=_�L�^_p_�[�ATB_�� $"��ipT��A_AWAY�C^
�GCP *�=���V_AL�@M��R�B�Y���*��H_�` �1���� , 
^7�6�Boo�f�P%M��Ij��\@��c�ONTIM��&*���fi
�$cMOTNEND��#dRECORD �1+"�er9�Q�O�Oq=6��R{� ��Hx��O�s (�:�L�������� �ʏ܏� ���$��� H���l�~������Ɵ 5��Y�� �2�D��� h�ן������¯ԯ� U�
�y����R�d�v� ���������?���� �*ϙ�N�9�Gτϧ` �^�ϼ���=������� (ߗϩ�^�p��ϔ�� ���9�K� ���!� H��l����ߢ��K� a���Y��}��D�V��h���RTOLER7ENC�TB�b�P�L���@CS_C�FG ,0k�gd�MC:\��L�%04d.CSVdi��Pc���cA +CH z�Poo�n�"W^m�c��RC_�OUT -�[�=`�o��SGN �.�Ur��#��05-JUN-�20 13:15� �Q25-M{AY�1:00 �af P�X���n �pa��m��PJP��{VERSIO�N �
V�2.0.11�kE�FLOGIC 1�/�[ 	tH�P��P��PROG_ENB�_r�WULS�g �V�_WRSTJN�`��Fr�TEMO_O�PT_SL ?	��Uac
 	Rg575�cO 74T)56U(7U'50y(t�"2U$tH�/z2$TO  >-�/{[V_�`EX�Gdu�3PATH A�
A\�/]?o?��kICT	aF�P�00g�Tdc�eg��1STBF_TTS�h�I�3U��Cda�6�@MAU� ��bMSW��1D0i�<�l� ��2�Z!�mO|3bO�O�O�O�O�O�O_tSBL__FAUL� 3�_|�cQGPMSK�^�bTDIA��4�=�d`��a1�234567890�Wc|6P�/�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o\SZpPf_ *��O R*�?%�PBhz� ������
���.�@�R�d�v�H|��U3MP4!Y )^���TRNBKS��ĀPM�E�5ЏY_TEM=P��È�3��D3�����UNI.��Y�N_BRK 5�����EMGDI_�STA%�W�NC�2_SCR 6G��_����͟ߟ�f ����0�B���~�e�17��;������¯�,R|�d�8G�� a�������N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶�0������@$<� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ��������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/� �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gO�/�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo�Oqo�o�o �o�o�o�o�o% 7I[m��� �����!�[oE� W�i�{�������ÏՏ �����/�A�S�e��w���������קETMODE 197��v� '��� �W�RROR_PROG %��%���X�'�TAB_LE  �A�𚯬���њRRSE�V_NUM ��?  ����)�_AUTO_ENB  #��j�w_NO� :��
��  *�*F��F��F��F����+E�_�q����HI�S�h���_AL�M 1;� �2��F�F�+�� �@�$�6�H�Zψ�_�.%�  �D�����ېTCP_VE/R !�!F�j��$EXTLOG_7REQ�������SIZ����TOL�  h�Dz����A ��_BWD��5��a�	�_DInO� <7���	�h��k�STEP�w߉�ې��OP_D�O��4�(�FAC�TORY_TUN���d��EATUROE =7�a���Handl�ingTool �7� DER �English �Dictiona�ry=�7 (RAA VisS� Master0��>�
TEa�nalog I/O7��>�p1
a�ut�o Softwa�re Updat�e�� "`��ma�tic Back�up;�d
!���ground� Edits�  �25LCa�mera��F�� w"Lo��ell���>�L, P��om�mj�sh�8�h6�00%�co����u�ct%���pane�6� DIFD�'�t�yle sele�ct�- `�Co�n��j�onitoir<�B�H��tr5�?Reliab�� ��(R-Diagnos���:�y��Dual Che�ck Safet�y UIF��En�hanced Rob Serv��q (V�U?ser Fr����T_iE�xt. oDIO ��fi��u Z�\=end �Err��L��  �pr�[r��C  �P���ENFCTN Menu��v����.fd� T�P Inp�fac��  
v�G��p�l�k Exc	 g�5t��High-wSpe Ski��_  Par\�H��~G mmunic��wons��\ap�ur� p���t\h�8��con�n��2� !D�Iwncr� strZ��i�<�M-6< KA�REL Cmd. L� ua���8~sRun-Ti4 Env=�(mqz �m�+��s��S/W�=�"y�Lic�ense��' a����ogBook7(Syo�m):���"MACRO�s,�/Offs%e��f���HG R����M1?�Mech�Stop Proyt��d 5
$�{MieShif���9�B6SD�Mix� ���7�y�Mod�e Switch���Mo����.& R�M�&��g' 6�5�ulti-Tp� ����Z�Pos���Regio�  �! 7Pr�t F�unb>�6iB/1��Num ��d�x�P`�312  Ad�ju:�/2HS�M7Z* oY�i8tastu1<�AD �RDMotN�socoveW� #���3�uest_ 867.�9oG �� �SNPX b����Z#Libr<V�;�rt IE,�� S$@�.�0�� ��s in VC�CM9��0�� `��!9�3��/I�� 710< TMILIB�MJ0,@� ��Acc����C/2�@�TPTX"+QTeln �Lq3�%�|(PCUne�xcept motn�� �0�0,	7�?\m72f�+�4�f�K  h6�4aVSP CSX�C9�@(P�U["3� 7RIN�We'g50,D��Rvr��	menS@� �Qi�P^ a0��3fG�rid�1play F O`�fp@���vVM-�@A(B2�01 f`2� O{RD|�scii��oload3�41%�ylJ�i�Guar�d$P�mP��k7�b]naPat�& 0N"�Cyc��0or�i���`iC00Data�@qug�c�3p[,`�3FRLOA�am�5<�3HMI� De�2(�1oc6�44�0PC�sePasswo�aA)qp��1p���{-+Pve�njCT���YELLOW BO�I� t�"ArcV0v�is���%���We{ld� cial�$_    �et�sOpA ;�41\\��5a 2��a��po0)@`@�aT1���5�0.2HT� @ xy��R:�82���`gp�P��xp�� 12�A�JPN ARCP�SU PR\A�T�Eh0OLwpSupg�fil5p�Q���^ l�cro�6 "AT�`�3ELdx�!���SSwpeetexn^$ J3�QSo��t� ssag�% 	T�eBP� ] !9M�Virt��39�V }h	`stdpn6����ro� SHAD~�pMOVE TF �MOS O � D�get_va�r fails ���ߐ  � D��E���� Hold �BustdCVIS� UPDATE �IR��CHMA �62�q�WELD}T�@S ) "��~�: R741-�kou
�b��m �BACKGROU�ND EDIT �Ò m41�0RE�PTCD CAN� CRASH F�RVRTO�Cra�.�s 2-D��r� �0r$FN�O NOT RE���RED � P�CVl�JO�P Q�UICK�OP �FLEN .pc��c���TIMQ�V3 ldm�PFP�LN: 燹 pl� 2���FMD D�EVICE AS�SERT WITg iC��sANġ�ACCESS M� �aŀo1Qu�i��<!�C"�US�BU@- t & rOemov��<�2� SMB NULAp�ܡ��FIXW��H�IN͑OL2�MO� OPTt�PPO�STwp��D��- �� �Add��adl. 	�io��$P:��Wu`.$ѠO��I�N��M��CP:f�ix CPMO-�046 issu5e�tJСO-|�2��130���SET� VARIABL�ESΐ�$O�3D �m�"view d�a`PWea�80b~. of FD ���u)��x OS-y1�p� h s v�D�5t��s ��lso �(� WAx���"3 CNT0 �T�S$Im�Z#c�a��PSPOT:�Wh�p��s�STY�܄At�pt�d?o GET_l���VMGR LO�0�REA�pC��M�`P�@ Y��0�EL�ECT��L��ING IMPR N����Rɰ̐sPRO�GRAM�RIP�E:STARTU�@AIN-��D��Q�ASCII�d�O�F L���!`PPT�TB: N��ML�Kdme�4��:�m�oW�all��R� �Nu�Qr� Angȅ��`d��thzo�n[� ch >`pܐ�r R2toun��H85@�iRCaylA�"Sign�0��pI,A�Thre�sh123�#.c��Hڰ : MS�G_P�єper �ࠡ��A�zerqo5P� A�  J�!fO�Imr � 2D�0�rc imm�`SgOME�s�ON�������0SREG:��^5� LB A�9�KANJIH�n�o��`c	��n 9dq�� -1o���INISITALIZATI��cwe��0= dr\ � f��aP���min�im90rec 1�lc0�:?!blem��ro��L�<3a �i� 09 ��b�d��w-� ݡ�0�w� uHQm@se�4SY�M��s���QЧ �090�Wlu� E�;BRe��jձ4�1����m ���Par��r@ G�Box f�o TME�ːR'WRI<���SY��k\k��F/�up��de-rela2Q�d��#5�betw�e�pIND��GigE snap��us5�spo Vn�TPD��DOs�~ġHANDL �`�Q�i�D��n�0 �f.v���Bop�erabil�` stmCQ��: H5@r�`l��L�
! ���m@ph�s U�IFL�PO>�FA�����ΑV7.��C[GT��pi�AsM��5pj�)@U��ine-RemarkO@�0 RM-�$ÔP�ATH SA̐L�OOS���v�`fi}g�GLA  �0d%���p��J� ki �q�ther�A� [Tr�`in�DW��4��2�7�� X�е�h��8`n;� C� R��:  6�d� y* it 35\k�wPay�a[2]_^�D1: g�s> �dowD2	SDIS�p�1�EMCHK �EXCE ֠�$M'F +  ��h�"��P��Վ�B0 c0e1Ȣ��me�� �c� !?��bP��� BUG��yB
:�@DŠPET��V0�0�T93X�XPAwNSI)�DIG��>��O  H5�P�CCRG ENC�CEMENT`�M�m�K 1A�H G?UNCHG OA�1�Tڐ����Sg\�d���10ORYL�EAK������L�C WRDN R���O�`j5`PO�S�PEްCG�V 7ont��VM�����W��@`GRI,@A�7��� �PMC gETH�0i�SUذ�>� H57�P0PENS!�N���ː� RE (i�RO�W<�³RMV ADD  II�=p���DC^ q�T3 A�LAӀ ��m��V�GN EARLY>���f n� ��衸E��ALAY7u�СPD�g�ˀH1SS8�OU#CH��D��Fh������PCDERROR�*PDE��� WRO���CURS�PٰI�p@N gҰ�?Q-�158Kwa���S�R �ġU3��\�aptp��@T�RF�@�R�\`�UB�U �`��#RB�0SY �RUNN���`10|�ఱBRKCT@q�ROq�Ԁ���CDA�X��Djj�EISS�Ucހ\��D��TS�I�aK�tXM�IP�SAFETY C�DECK "M6 ���dѤ�[`S U�)�8�4}P@QTWD��E��'QINV��D Z�O����a�sb_aBD�UAL@|�'QòFR��E�4l�6��P`?NDEX F�P�U,���SUF�rPk�Lb�ѳ�RRVO117 Ay�T��챤 ���FAL�BTP24�7���P?q�EHIG�PCC n��0�EoSNPX*PMM�QE ��)!SQ�"V���8T�bDC�BDETE�C��ds!Sˀ�BR�U/b63���s� 0C2"�t�s�'�!h� Z�T�7pS��"e���߆��,����߉ـ��0�
ա��ق�c�scr�ـ �dctrld.؁��$�fّ��!���qfـ*��878���-�% ��� rmґ�
�Q�R��78��RIـA�̑ (��~��Q.����ao�ـ\��a:P���a���I��ta 3 "K�:����<�#�o��t�p؁ "PLCF�"E!�ـ�plc�f���ـ-���maai�ـN���ovc���ـt�/�ـ����x��􁢐r674���Shape GeQnwـI��R,����ـT�іV� (5�ـ��II���� �`+��ـl���sga �4P� 4j�I�r)6ـŲ5=�5ѺI�n��ets6� " �PC���nga�GC�REѿ|�5��@�D�ATj���5ŝ�t.�!��5�a񯜳A�g�tpadb���Y�tput����������2ـ��5Ĺ���f��sl�q� 7�hexy��4����ώ2�keyy�ـ"�p1m������us9ߜ�gcـ����x+�H�a�j921��pl.Colly�����r�ВN��ڕr�3 ({�ـip����r��'���8�7=�7����tp�� "T�CLSj�|���cl�sk��D���s�kck���)�U����Ѱ�r�H���71a�-� KAREL U�se Sp�PFCTNj��7��a�a��� (��ѡ�� �ـ���ٹ�6�8=�8"�   �ـ 0�S�(V� �  lm� 6�9�9�~ F�)vmcwclmf�CLMl�0�`��60vet���cLM:����sp]�~�mc_mot����ـy���suX��60����joiT�J��_�logH��tr1c��ve%�� �����g�fin�der��Cent�er Fb!��M�5�20����g��  (�m)r,���fi ��1��a#z�� ��ـJ��$tq� "�FNDR����$e�tguid@�UID�ـ
?1��E7�q1nufl�60 �ـ>_z#ѯ 7A�x��(�2#���$fndr����c$���tcpS$]�CP �M� H�3ـ517��g�38�vC� gD�*Y=�F| Ց� ^ ����CtmgA4�P ��O�CG1ՑO7�Y��8�Etm �?�W�ـe�?�C�Rex��ے���Z��ڔXp�rm؁�_�D�_vars�_Z$M���V�h@����`�gG��ma|�w�Group�@�sk Excha�ng{@ـÖMAS�K H5�H5973 Ha�H5���`�6�`58�a9�a8��B�a4q2���b(�o#
k�/�غ`hp
8�0Y0/_цt�qTASKY_�r��pz�	h�Z�m@���������SDisplay�Im��v{Gـʑ8�OJq(P%���@xa���a�� ـ�lqvl "DQ#VL�t���q������Ϧ�y�����1av�rdq֏4ᩅsi1m���0��st��o���d���������v��0Z樁���"v�Ea�sy Norma�l Util(i�n4�|+11 J5C53��a�c���(���0��)�M�<�O�<� /k986TA8��#|�4�� "NOR�
`��1�_���|�su�� .������7���a!g�~y! menuu���g#M�����R57�7� 90 ̒J989��49�L�A0�(�ity�E�A�,`�P�m&��mh8��"8 2��܄����C�8_Sշ�n "MHMN�r%.Ը%� ��ͯ�s����i�Ը-at�Х_������֌ֶ��tm�?мz�1�����Q�2�Ͽ�z�3<zos�odst��
��mn�O��ens%u�Lm���hRaL��߃��huser!p�a����c~����Ը5�ɯ�����op�er���XԸdetbo`Ý~ ��L�UA��������dspweb���+�X�r��u<1��101W��הּ�2N�A�e�3!0A#0����4N�;2e�5��|����"��CalxN�0�O��Z� �0�O�$�S%j{�u���� 0S��}���ump��\b�bk968�!68�!��b�eq969B�9�%��F0b��? "BBOX�ۍ>�sched����setu~Xk��� ffH)�0��eq)��0�col(�1bxc��8�li�Љ�aI����W!i�e@m�rof$T�P EB!TA&@ry�|M427�*l!(T\�Q!RecX"H
�q�z�?$it%�?#сk7971�!71�{�F��$parecjo���A��?'����X�rail�@nag�e��~@]��D2E� �[0 (?:H͒V|x@@1ipMa���3�p�!�4�"4�u��3pa�xrmr "XRaM$��3�rf����ß1�1ꫝ0�yturbsp'G#��^@� �015: ��625t/~A��\BH�'ZD iy!:k�E�6�"A���H� �7��P�.��E!pd "TS�PD�}�T�GtsglD��kY��O�CiC�sRct%���Hvr�vQ���K�P,��A  q#-a�21�Y@AAgVM �r-b0 ��fdE`TUP h�im (J5�45 l) �i`6�16 V2VC�AM .CLwIO Y10k �5W` (F�`MS�C ���bPs��STYL�Sua28y kr�`NRE I��`SCHgRp�DCSU tps�h ORSR� �ua04��EIOCW`\fx��`542 LEX="�`ESET��ia,y`0shi`7y`"R?MASK�b�7o�-`OCO[�x��a7p3Sv q`t7p02kv6U`xv39_v�x�LCHRvOPLG��w03;uMHCR�3MpC�`YaP`�p66�.fia54; #��MpDSW�`588��ip1�a37 8/8 (Dr0c�5r94���r7 qj5r�5�5r^v�p5�"9PRST VR�FRDMC�Sx�a��-`930 �>�`NBA  g1�`HLB 3 (�a{SM�� Con�`�SPVC Lia2�0�#-`TCP a�ram\TM�IL r�PAC�C�TPTX �p��`TELN 96��0�r9/uUECK��1r�`UFRM setL�aOR ���`IPLKeCSX�C�pj�qCVVF� l F7�HTTP strbZ0zcp�CGy�8�AI�GUI�p7 ��PG�S Tool�`H?863 dj��q�M�Oq3
vJ684c�\$���sق��s'�1ےs�a96� TFADȑ65�1�Cq53 � oo�b1�44r-�k��r9�VAT��JO775 �R�6u�AWSMے�`CT�OP �q�`olld��a80;!diy�sXYY�0 e���i`885 '��`LP�`u"�`� 7H�`�LCMKP��pTS�S J%�
�W�CPE \dis�`�FVRC m��N}L�U002 
�{en%�6 65JrZ'�7[�U0�po��Ƞ�K���t� I�4 �URI�5�&�U02�2 nse�{�3� APFI�`{�4b�2�`-���alOP���1C�33O�͐t�ptsD`U040&g�43�ٲ4�۰j� "sw%�1`b�	�4�C	�5 ��w�x�57�eU061t��S�6ұrob9�15g�i��68����$!!��7�w�7�Ё�|%���"rkey��	3w��4?ǽ���T����8'�089�U#09���P��9:����2 &�l �9&�l2��9B�VrU15�P�NM� slA �3#H�}���1q�0v4ӽ7��108 	�eDэphc ��s�1�q�4+�1����A�5J/�tx�1����1]p!u�Qѡ�t�1������`��3����6��1�!p �`�о�- W�8�147 ase� C�U`sB�1 �82��1�4�8� (Wai��599 ��aU166�W��1�W�4� j U�6$�#U�7�3U�8�3�ȱ��B��1{��2 �act���6 "M#CR@�ِ4�1�������967ǑU1S93�3��6��2Y�dsP��2A��21���as�F���<�28-���E�2 wF���Q55�(��� ��cر5)�w���q��p����qf��L��$������q4d��2g�8q��8�51�""]�}�q��"< b������B]� � f�; `�̑ � ?8 16 (ݰ �BA��AAҰ�]���g :�!��`8 bbfo=� t� �j�� 7 \�� ]�� �2 �k_kv��74 0&!����W0H5���57&�579 h� L82 %"�\�4 3��5���5��1��59s4 U219 7,�-�6�p��6i�\t�chH6ur% �4>S3� 90� h��&�\j670��q���r!tD��4��&�t�sMg�lc�S�FrE�H��#F�����hk$�� sC� � ��"F�L��dflr��� �� ���fu!l%Z�gvPva���� sA����"D��3|��!creex�� �!�%�!�%�,���6�j6�s�!prs.�!�%�!5�hA�x�P 5�fsgn���/�/�,at<D�AD����qs`R svs�ch`@Q!Servwo S�!uleoCnA5SVS�!44�0��F��1 (�0A/ched�0,1�EA၍�� �2Q��0@��^�r0�U)1BBc��+� %P5)Q1�V�-#�3�1css "ACS�WVY88"gA@�`8!�/�0��@e���#M��C�3�tor�chm�0�- T�QMa�1�1M%'�9� J5lA598 *א1�!7)P8<P(1�̢A�ء%R1Qte,�!)E A5E`AS�v�� mLC6AR]C_� 1�4qc� �V�Ht!tc��A耥Q�4��R �F1 7T!2�S�EPBPQf-!�RtmkQ!p@60X��/�PRC8S�Q#�S�) P�2a96xAn`X�D.<bH5�1�U�}E� T�Qf#` aQ!<���F!�T!!�a4�3FcRO�Ttm�R!av`58�_�WP��MA$q�E88��>rp�in_��(�o�@e`AcB�rr��)u�!�U�etd�ѧ�U�Qovet�o�#$,�S�mmonitr42�=�Q�cF�st,"M_va�P`47M��V�0�! 5�8q���ameQ!Ɂ�rol�A��43�$Q0  Sp��1�0�1$P25�AKR  ��� 0S��(V�Ɂ)xj818\nl`mD��zN���r�MPTP"��O��qmocol �]/
�Y1�4Xa�@䁘�2�0i�53(1��T/ouch�!sؠ�2%qD2J5 !IU�٠��= b�0n��A�� ]�vP���z�EOWJ�th��Kwc���{��etth8!TH�SRXâm�t�o? "PGIOsRd�'z�wk� "WK�1�aL&MH�PH5�4�5�Q5�o��m`A��q@7z@6���1�8�a�PMor��tsn�@T�A�o�c���P"�����m�uA��T��p���T?��|�m4�TM�!2�5 4�>����m9�w�f�h�S�3G�qor�3���"641���8���Q!A�,HE!pR�U <�m�Re�h-g? "SVGN_��(�copy "CO�TA��U(��r#j0 "FSG��_�eh�j�f�@wA�SWwj|RbY=sgatu����!�;B�tp�AT�PD7��9 a790s����sg8!���GAT&o<Rc9  �Ħ�1�@t2`%1�&��1�bpv �1��&�1��B �1�8 6�1�chr��1�|v�1�sm��1�v����gtdmen�ps1�(v0!1��mkpdt�r1��]A1��pd��1�$&��1��mvbkup�.1��6�A��mk3un��G�pr���Gmkl1�e�P�s1��ni��0&1�ldv9r���glg�t��1��&���#�auth�.p�&��1�����) sud�1�7@� 1�G�1��\1�g b2�p�w 1�x6O�Ł4� 1��Ђ   946�"1����1�t\p�aic\p4k9471�wc��1��ictas-�Mpa�cck0m	8�	gen!1�I wl��Q� �stfq��q�wb���������vri/�4�^���B1�D��Pflo�w�@��Ac0ow�3<R50?���Q�TR�  (A0e T�0)B�Ԗ�cud!�0w�1��z�ac�$0�46 a� =�f�+p�aRa���!1�355Ţ1�F�ѡ�)a%|��;:afcald�� �&�0����%�f�m:�"�#�4�`��'a`"�3U���$��B1�! trac�k���@aine/Rail TrP̎�{(69�/�@ (L !iEYB�ʔ_ VB!Bu��a YB38P�48'7�	�F2���4��/�C�B1�3bŢ3�/�IUal��1�NT����VA��zQ�in�p�?0HVaen0�?DXWApuA�8�YqBzQtstd�0 U�@1GW ��]�j�VD����E&��VH@���o�peners^CO�`�ADev/w'~6�F8��񭁶��bA��aes�#1�]�ג��d����m�d1�k)9�@7�6��#1���/b�epaop`aO�PN�Wj�`��Krc#el}?�Exg���Y8`5Dv��tscx?tб�a�s FuvrCop /�Dw�nDh ��bAr5��QB�g�d�k�j!�� Pump v$Aᛑ�/�1�a;��M��T�q�i����t4U�1� 0�S��O \mh/plug�gr7G�h���u|bZ#��io�h#C{p��v(�ALI�O1�1�@7��93�Q51�91�����]4�� ST�
R��t�J989��/RL�SE�g1�@Cd�(M�1�/O�'�Q�)�D��G1 zq�H1�55'?��zq�tcwmio��MIO��$�tc�q"CL�01�UQcP�|�iEo��u~0%�l9� zp��v�1o���bQ�tzt����dtz�5I$��V%�rh#Inste�Q�� Co~PIo�qvRP1�hd�B554 (l�oBv��,�Q�H��Tcipc��oo�ڱp5�A�(
@��������"7`����aڰd�QCD �W�	����8��ڱ�rGcnd�_׳1p�a�ײ������Sb��a��O�2kz<�rpcrt�ᱯ�pٱdEc��S d��\���u�E!߳vr2k�pE A�-�x�_B�\"� choO�l"u�C��Y 1খ630 @ᗷ�@�� �ӿ�q�X�ԑ�GTX�? ��>�1chp "��XOh:�3�&�"5x!E��\p3 ���P��j�d 11�$h��Plo���ұ�c!h��3��s1��a�01���#Ar�� �0� !oCB��spq[`Jm:�k�7�)�vr�������a!X%-J�FR�AJ�Watpqrn�ev'�����fQ��D5��`��KrboT , �$��PG�[z!�sm�ICSP\Q�QP5y��!QP���j�H51�z�93QP7y�6���������5��R�6QP���NPR�`(�P@aam S`u��b��ĉa4tppr�g�p�B�	�Z�qratk932(q v輏�sc "iC8��~�atpr�_��qqz�;F�LGds�blflt{�ёs�able Fau`��CPav�aQ��~`aDSB (Dt$�t�d�A����QPh"@�E1��`f$*��3[S�� A�"tdj  "`PaV�Ohf$�1sbj!��1�"\:1gc��.��f%�du�550^CA�djust Po'int�b��J/��-��0�4�a昐A��j��O�N0\sg�4x��w�1\ada��O"ADJ�M�j0��etsham�SH�AP0���XDjpo  �e��G�a��UGQPG'(.��1:�k@ab5�J��KAR`�iagn/osti��!�a��66 J�C��a=P�(QL�Q&T�o�fkrldeP@���	  ��SQ��)�3/ρ[ypp��DBG2t�!O �U�Rѯ#��V��F( �шS7��Q�i�p{�M�ipper Op��Pq�����78 (MH G w�1Rlbk_�fTcBQ���0&�d038<B8�t��E��c�9_9�t��Tc��k����8 $q�SdrnpVǁ� �Qd�Ő6Tea�=����r Mat.Handlv �an`W�� MPLGv�A_�p�q(�sє�f����g ��b��a���f�� ����>@$w���� Dw��EI d���uu��m���fhnd �"F��  ��)���#� ��p���>��(Pa�0To�@�$V�!!�3#p��a�>��{�Q�k925B��26�q�3�{�p���2	ş�y���gse>0GS�qďėPR���T���a���t�p����{�dmon0_�q�Ŗ�ans���vr��{�=�����ͪX�<y��wsl� � pen��D��Y�WA��823X�Q
� G�0!'�&P��8QqI�Q�GQ �\sl ��!q��v����������֐�_�`����"S�EDGiOٳaQ�tdg�@T�AF8�F�� �BN���ÑQm�7���ڱA��g;Ж�Q���8��q�S�ileg�y�e���ϟ�9�F'QQ�<LaQQj517So�3-[JV�?�'�#4BA�49GA�WL�aw {�no�Qfԫo�H17D�#a������0t�  �>��LANG j�A5��5�5� gad5��C5�,TC5�jp .5�ce���5�ib=�5��#5���pa5��C5�W�~��j539.f5��]QRu5� Env�
5�5S��K�3y ��J9$5�.� ��;��G5�2D2�5�JS��p(K}�n-Tim��"���"¡�3H􅓹���\k}l5�UTIL"������r "QMG���,q5�C5��1 �"5�ړ5�s5�\kcmn��+��r5����utM�_�lre3ad���ex����"��\��l$"��1a35�rt[! -5� tuva��`_��5� �`CV����\�p ���Bp9t�box��_qcyscs}kRBTv�veriOP�TNv��l��e`��K���hg/>�agp.v1$�"�1$ptlit/DPND�BPm$d>n#te\cym$8$xo"��#mnu3�/�/�/�.5�/�/m$���UPDT it�e��.3 swtox95]�-4oolBD5 wb95��-4FR-4Y�� /2grd�-4��-4�b-4��w-4B-4.3 ��-4�-4'�-4�.3�B0l� /2bx "`�5�Q5I.3tl�7`��AE�#/2r l\�6��@O�-4 :4CoElD5eMa-4+�C�5�K�-4W�Q5ml�-4Chang95}�95�qQ5rcmdE�b�OZ��`6�5,r�7�6��70�5&r_+]22=_O]!2� c_u_3U4<_N^�57�_�_1UCCF�M�Ey��_accdau59#�6cAEX`� /2|�Da��4|aO/Jm�a�5�-4@�4�a AOSJ	Q�e�o�o�Y��-4��ZDQ-4sQk��?�@rtet�q�-4\$�3�q�eunc�.-4��4�q�5su�b�5��5E�q�5cce�@oRf^opm4E�o�fv�7�o�eT �c �o�nt$
Pte;�q �@�f\��k��6;��-4Ѓ -4�K�D��zh!-4xmoQv�b�q�et����f�"�tgeobd�t.���ƥ�etu � ɐ��ɐ��tɐٓ�xߟ�z��va�r'��xy&��pclJ�cɐ��ɐ��eɐgripsu����uti�����infpo��ܯ�B��ɐ������\�����ɐ�Ʊ�8�p��n ��ɐ%�ɐZ�mT���0ɐԶ��\�ogġ��p��%�p�\�palp�����s����ɐݵ���Ŵ����p�p����p�kagd�%�7�lclayY�k�A�ɐ��Adɐ5�p�������B��|�|�������q�����rdmͿ��r#inT�-�?�sO�Q߈c�̿޼s���ߧ�t�v�ߧ�h���s�tn[`��tX01�ɐ)�Dɐ� �Tu!l4�q��g�26Ϥ��upd����vr����נ1}�3�נ�ᜣϵ�il3C�U�l4����T�5e�w�s �ߘ�֠�߻�wcmx�(��xfer�~��tlk2pp���conv�朗ccnvݑ��5�ag, y�lct���n�yp��nit0���d���(��  ��ɐ 0S�(gV�U9al �#pm�Wse��2� ���V�C��(�z�@��A�0�|�m��`��&$��޷'#ro��@T/f(&���p1�mI� �,��$�+���/ �)G�?�+�� �L�ɰm ∡P?b6D�4 rg�������� ���?�9�� O�7�� ����>�/�T� a�8/�C�����E��b,֡)?�*��nq?_9�l�-!H�� � �HA |�p��QU1 p! �O���P ��S i	�Q�R@t�`�  ?���ɐ8� ��M�.Oreg.�ԃnO�o99� �� ���$�FEAT_IND�EX  �S �_��P�5`�ILECOMP �>���ba�Pa�RUcSETUP2 ?be�lb�  N� �aUc_AP2B�CK 1@bi � �)�R�o�o # %�o�o�Pe`�o )oe�oU�oy� �>�b�	��-� �Q�c��������� L��p�����;�ʏ _����$���H�ݟ �~����7�I�؟m� ���� ���ǯV��z� �!���E�ԯi�{�
� ��.�ÿտd������ ��*�S��w�ϛϭ� <���`���ߖ�+ߺ� O�a��υ�ߩ�8߶� ��n���'�9���]� �߁��"��F����� |����5���B�k��� �������T���x� ��C��gy��,�P��qi�`P�o 2�`*.cVR�H� *K�q�w��2PC���� FR6:D���/�T@` @/R/�=/|,C`/�/�*.F5�/�	��/ <�/$?�+STM D2M?X.��E?�=� iPe�ndant Pa'nel�?�+Hz?�?�j7�?�??-O�*GIF7OaOl5MO
OO�O�*JPG�O�Ol5�O��O�O5_�
ARGNAME.DT?_��o0\S__� ��T�_@_	PANE3L1�_�_%o0�_o�?�?�_2orog `oo/o�o�Z3�o�o@g�o�o�oH�Z4�zgh%7�KUT�PEINS.XML�o_:\���q�Custom T?oolbar(���PASSWOR�D��FRS:�\k�*� %Pa�ssword Config����� ���+��O�ޏs��� ���8�͟ߟn���� '���ȟ]�쟁��z� ��F�ۯj������5� įY�k��������B� T��x�Ϝ��C�ҿ g����ϝ�,���P��� �φ�ߪ�?�����u� ߙ�(ߒ���^��߂� �)��M���q��� ��6���Z�l����%� ���[��������� D���h�����3�� W������@� �v�/A�e ���*�N�r �/�=/�6/s// �/&/�/�/\/�/�/? '?�/K?�/o?�/?�? 4?�?X?�?�?�?#O�? GOYO�?}OO�O�OBO �OfO�O�O�O1_�OU_ �ON_�__�_>_�_�_ t_	o�_-o?o�_co�_ �oo(o�oLo�opo�o �o;�o_q � $��Z�~�� �I��m��f���2� ǏV������!���E� W��{�
���.�@�՟ d������/���S�� w������<�ѯ�Ơ��$FILE_D�GBCK 1@���ʠ��� ( �)
�SUMMARY.�DG篓�MD:��[���Dia�g Summar�y\�i�
CONSLOGQ�4�F���߿�n�Consol�e log�h��G�MEMCHEC�Kտ��J�c��M�emory Da�tad�l�� {)}O�HADOWY��>�P���t�Sha�dow Chan�ges��£-�?�)	FTPҿ?����C�n���mme?nt TBDl�l��0<�)ETHERNETaߑ�"������n�Ethe�rnet ��fi�guration���s�V�DCSVR�F`�F�X�q�t�%�6� verif�y allt�£1�p�1�DIFF�i�O�a���u�%��diff���"��6�1������{� ������	9�CHGDE�W�i���u�!�&��9�2������� ������GDM_qu�8.9FY3���� ����GDUgy/u��6/�UPDA�TES.U ;/���FRS:\S/�-�o�Updates� List�/��P�SRBWLD.C	M�/��"�/�/���PS_ROBOWEL��g�\?n?���? ���?�?W?�?{?O�? 	OFO�?jO�?{O�O/O �OSO�O�O�O_�OB_ T_�Ox__�_+_�_�_ a_�_�_o,o�_Po�_ to�oo�o9o�o�ooo �o(�o!^�o� ��G�k �� �6��Z�l����� ��C����y����� D�ӏh�������-� Q���������@�ϟ 9�v����)���Я_� �����*���N�ݯr� �����7�̿[�ſ� ��&ϵ�7�\�뿀�� �϶�E���i���ߟ� 4���X���Qߎ�߲� A�����w���0�B� ��f��ߊ��+���O� ��s������>���O��t�������$FI�LE_ PR� �����������MDON�LY 1@���� 
 �5�Y� 0}�=f/��� �O�s�> �bt�'�K ���/�:/L/� p/��/�/5/�/Y/�/  ?�/$?�/H?�/U?~? ?�?1?�?�?g?�?�?  O2O�?VO�?zO�OO��O?O�OcO�O
_��VISBCK������*.VD_[_�@�FR:\F_�^��@Vision� VD file �_�O�_�_�Oo�O)o �_:o_o�_�oo�o�o Ho�olo�o�o7�o [m(� �D� �z��3�E��i� ����.�ÏR���� �����A�ЏR�w�� ��*���џ`������𨟺�O���MR_G�RP 1A���L4�C4  B�9�	 �񝯯�����*u����RHB ��2� ��� ��� ���ݥ������ ���ި%�ߤA�5����_�J�KsӦI���HhV�T���}R�R�P����M���q� �F�U<Hp��G,*;��h�;r��@N�-ޝ�@�2���2���E�� F@� %5U1ŝ�J���NJk�H�9�Hu��F!��IP�s���?@�u�ÿ9�<�9�89�6C'6<,6\b�������������� ��A9�A� ?�M��r�ߖ߁ߺ����  >o"A�\a@��@���߳����8� #�\�G��k���������4�BH9� ��8�����>�P��`�
��P�X�P��k`�w�����B񤓠��M�@�33���������UU�U!U<�	>u.�?!����k����=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:��7p��D�@ D��� C�@�UC���Ώ�'���� ���-�/�C/�#/ 1��/Y�/�/�/�/�/ �/�/0??T???x?c? �?�?�?�?�?�?�?O O>O)ObOMO;�N�P� ^O�OZO�O�O_�O+_ _(_a_L_�_p_�_�_ �_�_�_o�_'ooKo Xi�Xo~o�o�oi��o �o=o�o�oBT ;xc����� ����>�)�b�M� ��q���������ˏ� ��7�/{/%/7/�� [/��/ܟ�� ��$� �H�3�X�~�i����� Ư���կ����D� /�h�S���w������O 㿩�
ϥ�.��R�=� v�a�sϬϗ��ϻ��� ����(�N�9�r�]� ��]o�������߷o� {�$�J�5�n�U��y� ������������4� �D�j�U���y����� ����������0T �-��Q��u���� ��ϟ5GP;t _������� //:/%/^/I/�/m/ /�/�/�/�/ ?ǿ!? �?Z?E?~?i?�?�? �?�?�?�?�? OODO /OhOSO�OwO�O�O�O �O��
__._@_�d_ �O�_s_�_�_�_�_�_ o�_o<o'o`oKo�o oo�o�o�o�o�o�o &J5nYk� k}�����1� �U����y���ď ���ӏ���0��@� f�Q���u�����ҟ�� ����,��P�?q� ;?��[���ί���ݯ ��:�%�^�I�[��� �����ܿǿ ��� 6��OZ�l�~�E_Oϴ� ����������2�� V�A�z�e�w߰ߛ��� ��������,�R�=� v�a��������� ��'�I�K��7�9� ?���o��������� ��8#\G�k� ������" F1jUg�g�� ����/�/B/-/ f/Q/�/u/�/�/�/�/ �/?�/,??P?;?t? �?MϪ?�?�?���?O k?(OOLO3O\O�OiO �O�O�O�O�O�O�O$_ _H_3_l_W_�_{_�_ �_�_�_�_o�_2oDo �eo/����oe��o�� �o��
%o.R= vas����� ���(�N�9�r�]� ��������ޏɏ�� ׏8�ӏ\�G���k��� ����ڟş���"�� F�1�C�|�g�����į �?ԯ�����?B��� ;�x�c�������ҿ�� �����>�)�b�M� _Ϙσϼϧ������ ���:�%�^�I߂�Io [o��o�ߣo�o��o 3��oZ�u�~�i��� ��������� ��D� /�h�S���w������� ����
��.���� '�s����� �*N9r] �������/ ۯ8/J/\/n/5��/� �/�/�/�/�/?�/ ? F?1?j?U?�?y?�?�? �?�?�?O�?0OOTO ?OxOcO�O�O�O�O����$FNO �����A��
F0Q �P T�1 D|����@RM_CHK�TYP  �@�\���@��@�Q{OMP_MIN"P����NP�  �X�@SSB_C�FG B�E ��{_���rS�_�_�ETP_D�EF_OW  ��-R�XIRCO�M!P�_�$GENOVRD_DOCVs���lTHRCV� dedd_EN�B�_ `RAV�C_GRP 1CdW�Q X�O�o�O �o�o�o�o�o& J1nUg��� ����"�	�F�X� ?�|�c�������֏�������0�bROUrp`I�HQP������R��8�?T쀟3�|�������  Dڟl��6�@@�B����p��o�4�g`SMTmcJtm蕗������A�HOSTC]R1K�O�pP�a� 5M�����0�  27.0G�=10�  e'�t� ��������b�ۿ�����4�˿ų	ano?nymous8�fπxϊϜϨ����л� ��%�'��[�0�B�T� f�x�ǿ�߮������� ��E��,�>�P�b�� �������������� �(�:���^�p����� ��������� $ s�������� ����K� 2D Vh�������� �5GYkm7/� v/�/�/�/�/�/�/ ??*?M/��r?�? �?�?�	//-/OA? c/8OJO\OnO�O�/�O �O�O�O�OOM?_?4_ F_X_j_�?_�?�?�_ _%O�_oo0oBo�O foxo�o�o�o�__!_ �o,>�_�_�_ ��o��_���� So(�:�L�^�p��� �o��ʏ܏� �u�١�ENT 1LO�� P!��E�  A�3�p�_���W��� {�ܟ���ß�6��� Z��~�A���e�Ư�� ������ ��D��h� +�=���a�¿��濩� 
�Ϳ�@�/�d�'ψ� KϬ�oϸϓ������ *���N��r�5ߖ�Y߀k��ߏ��߳����?QUICC0!����p�3�1q�M�_����3�2�����!?ROUTER������`�!PCJO�Ga�<�!19�2.168.0.�10:��NAME� !"�!RO�BOT���S_C�FG 1K"� ��Aut�o-starte�d`tFTPk H���s���� ��$�'9\ J������Jv !3E/Y{1/b/ t/�/�/g�/�/�/�/ ?'/�/:?L?^?p?�? �?Qcu�?? OO/ $O6OHOZO)?~O�O�O �O�O�?kO�O_ _2_ D_V_�?�?�?�_�O�_ O�_�_
oo�O�_Ro dovo�o�_�o?o�o�o �og_y_�_1�o ��_������o �&�8�J�mn���� ����ȏڏ);M_ a�F��j�|������� ��֟����/�ɟß T�f�x��������� !�#��W�,�>�P�b� t�C�������ο�� ���(�:�L�^ϭ��� ѯ������� �� $�6��Z�l�~ߐߢ� ��G�������� ����T_ERR M���.�>�PDUSI�Z   �^����U�>n�WRD �?���  �guest \��������������SCDMNGRPw 2NX�����p��\�K�M� 	P01.�14 8��  � y��}�B    ;����� ����������������������~��\��������|���  i�  �  
�ډ�ҕ�����+��������
����l��.�
��"��luop 
�dy�������&�_G�ROU8�OM� e�	0�p�07�	QUPD  �ŲU��!TY��M�@�TTP_A�UTH 1PM�� <!iPen'dan�������!KAREL�:*���KC����VISION SET� ://���Q/?/i/ ��/{/�/�/�/�/�/�"?�/>YCTRL� QM�P�v5��
���FFF9E�3.?��FRS:DEFAULT�<�FANUC �Web Server�:
Y���A<�OO*O<ONO`O<�W�R_CONFIGw R<� �?�>�IDL_CPU�_PC�0��B�ܩ��@�BH�EMI�N�L���DGNR_�IOG�|��S�@N�PT_SIM_D�OV[TPMO_DNTOLV 3]_PRTY)X�B�DOLNK 1SM����_�_�_�_�_�_|o|RMASTEP�&|R_O_CFG�"o4iUODEo6bC�YCLEdo4d�0_?ASG 1T<���
 o�o�o�o�o !3EWi{�p��k�bNUM{��Q��08`IPCH��o58`RTRY_�CN�0
RQ�6bSC�RN>{�Q�U� 6ba`?bUM��p�����$J23_D_SP_EN� M���ᆀOBPROC���LUMiJOG�1�V�@Q�8��?��{?ŃP�OSRE��VKANJI_`d�
_H�$�V�W�L}6h�1�C�CL_L�@�r��H�EYLOGGI�NB`���Q�PL�ANGUAGE Y�6�B�4 ��>�LGW�Xf?�ҧ����x% ���?�Z�@���'0��`$��>MC:\RSCH\00\�?��N_DISP YM�Ĩ�|�z�<�gLOCGR�BDz�D�A�OGBOOK Z�kR�P�T�X��B�T�f�x�����������v6	�<��⸥����_BUFF 1%[�]� I�2��H� S�h�d�n��ϒϿ϶� ��������+�"�4�a� X�j�|ߎ߻߲��������ˀDCS ]>� =��;����C��5Y�k�}���I�O 1^�k t��� ��������� � �2�D�X�h�z��� ������������
@0@Rdx��EP/TM  GdR2� ���0BT fx��������//,/>/)Ĩ S�EV:����TYP���/�/�/ ͆-�RS�0��*�2�F�L 1_��@�� 9�9?K?]?o?�?�?�?��/TPѐ��">ݭNGNAM��p��tU�UPS��GI����E�A_LO{AD��G %��{%��_MOV[��aO�DMAXUALRM�w��x{@AdQD:�<��C��y@C��`��Oj�lM�@̀Ҁ]a�k �X�	�!+�p+e���OΤ ,RX_C_U_�_7�|_�_ �_�_�_�_oo;o&o _oqoTo�o�o�o�o�o �o�o�o7I,m X�t����� �!��E�0�i�L�^� ����Ï�����܏� �A�$�6�w�b����� ��џ���������� O�:�s�^�������ͯ ���ԯ�'��K�6��o���d�����ɿ�GD�_LDXDISA��0���MEMO_{AP�0E ?a+
 � ѹ%�7πI�[�m�ϑϣ�y@I�SC 1ba+ �����'T,���
ߺ� C�.�g�Nߋߝ�߬� ������	���?��� N�"�������� b������;�&�_�F� �������x����� ��7��F� |���Z��� 3W>{���p���/��_M?STR ca-%�SCD 1d͠ �m/��/|/�/�/�/ �/�/?�/3??W?B? {?f?�?�?�?�?�?�? �?OOAO,O>OwObO �O�O�O�O�O�O�O_ _=_(_a_L_�_p_�_ �_�_�_�_o�_'oo Ko6o[o�olo�o�o�o �o�o�o�oG2 kV�z���� ���1��U�@�y��/MKCFG �e--��<"LTA�RM_��f��� v�����>�METPU�n����5)NDSP_CMNT������#�&  g-.a��v���y���#�POS�CF/�:�PRP�M.� �PSTOL� 1h��4@��<#�
��t����� ����/�q�S�e��� ����ݯ��ѯ�����I�+�=��i�#�SI�NG_CHK  �ǟ$MODAQ�Ӄi��a�����DE�V 	K*	M�C:�HSIZE��--ȹ�TASK� %K*%$12�3456789 �V�hŷ�TRIG �1jK+ lK%%�a���  �����όM#8�YP#���5$���EM_INF �1kڇ �`)AT&F�V0E0��a�)�I�E0V1&A3�&B1&D2&S0&C1S0=P�)ATZaߵߜԁH����p���	��A��9���]�D���  G߸�k�}ߏߡ���� 6�m�Z�l���K��� ��������� ���� ��hs�-�����} ����@R v);M_��� +/*/�N/	/r/�/ k/�/[m�/��� &?8?�\?�/�?;?E/ �?q?�?�?�?O�/4O �/�/??�OA?�O�O �?�O�?_�O_B_)_�f_��ONITOR�J�G ?��   �	EXEC1Tp��R2�X3�X4�XQ5�Xy��V7�X8�X9p��R0Bd�Rd �Rd�Rd�Rd�Rd �Rd�RdbdbcU2h2'h23h2?hU2Kh2Wh2ch2ohU2{h2�h3h3'h�3�R��R_GRP_SV 1��>ї��(q�������Yp�?�=
�҅?�OȽ�3f��@�_DR&����PL_NAME� !��p�!�Default� Persona�lity (from FD) ���RR2-q 1m)deX)dh��q7�X dv� ��$� 6�H�Z�l�~������� Ə؏���� �2�D�V�h�t�2������� Ο�����(�:���<��d�v����������Я�����*��R�,r 1r�yհ\���, �����~f� @D�  z�?���f�?�������A'�6z�ܿ��;��	l��	 �xJ԰�����˰ ��< ��� ���IpK�K� ��K=*�J����J���J�V尻�"�ɱT��:�L�Ip@j��@T;fb��f��n���%�4��=�N?����I��g���a������*��*  ´ [ ��P�>��������n�?z����n���Jm���� 
�ғ�%Ӱ�Ī�9��� �`_�  P}pQ}p}�}p|  �r��/׈�+�	'� �� ��I� ��  ��J�:��È��È=̣����6Ç�	�В�I  �n �@
�+�l�$��l����9�A�7�N�p|� � '��_���@2?��@���f£��@��C��C�pC��@ C��C��Cz��o�
�A�q���P @�*��
0�B�p*�A��2���`�o�R�n�Dz��q��߁��������2��( ?�� -�����������o� �䥵!�o�M� �?�ff ��/A>�� ��v��7�a��
>��  	P��2�(o��e������ڳڴD�?��o�x"Ip<
6�b<߈;܍��<�ê<� <�&�KN�A둳��nO�?f7ff?�?&�3��@�.��J<?�`�M�� ��.ɂ�����lƴ a2//V/A/z/e/�/��/�/�/�/�/8�F�p�/4?�/X?�y?��K?�?��E�� �E��G+� F���?�?�?O'OO�KO6OoO.�BL��B �_0���OUO[��O cO_o?5_�?\_�O�_�_�_�_U
�h��<V�W>�r_o�n_/oo,oeo�GA��d;���CRo�oNoD������o�o%�5yķD��8C|�spCH5"Z�d��y��a�q@I�~N�'�3A�A�A�R1AO�^??�$�?��;���±
=ç>�����3�W
=�#���{e���n�@�����{����<��~�(�B�u�����=B0�������	��H��F�G���G���H�U`E���C�+����I#�I���HD�F���E��RC�j=�z�
I��@�H�!H�( E<YD09 ڏ�׏���4��X� C�|�g�y�����֟�� ����	�B�T�?�x� c����������ϯ� ��>�)�b�M���q� �������˿��(� �L�7�Iς�mϦϑ� �ϵ������$��H� 3�l�Wߐ�{ߴߟ߱� �������2��V�A� z��w��������@�����R��q(�qg��������e��v����a�3�8������a4�Mgs������IB�+���a���{�&&	fT�Px���eP�P��A�O	\���*<��R^p��X���  ��� �*//N/</r/�)@�O� ��/�/�%�Q��/�/�/??'?9?  N?l/�?�?�?�?��?�2 F�$N�Gb���A��@Xa�`rqC��C@�o�TO� q�{OF� �Dz@�� F�P D��]O�O�I�cO�O�O__1_~�c?���@@8Z�^4� � �:� �n
 8_�_ �_�_�_�_�_oo+o�=oOoaoso�o�zuQ ������1���$MSKCFMA�P  R5� `6uQqQ�n��cONREL  ���a� �bE�XCFENBw
8�c�e qFNC't�JOGOVLIM�wdprd�bKE�Ywsu�bRU�Nc|su�bSFSPDTY�p)vu��cSIGNtTO1MOTeq�b�_CE_GRP [1sR5�c\:� I�2�m���Di���a� Ώ��Ï���(�ߏ� ^������K���o�ܟ ��ɟ�H���l� ~�e���Y�Ưد������F�`TCOM_C_FG 1t�m�V�8�J�\�
�_AR�C_$r�2yUA�P_CPL��6tN�OCHECK ?=�k �׸ տ�����/�A�S� e�wωϛϭϿ�������kNO_WAITc_L�w�e�NT ��u�kw[5�_E�RR!�2v�i��� ߠ߲߾��c���ߴ�T_MO�c�wj�, �V��3���PARAM:d�x�k�tV#ﰅ��=?�� =@3�45678901 ������������+��U�g�C�����y��������t���UM_RSPACE�o�lV>H�$ODR�DSP��v2xOF�FSET_CAR9T��yDIS�y�PEN_FILE� jq^�+�v�OPT?ION_IO�Y�PWORK y'�5s x�
fR�`"�2��2�	 �	2���[ RG_DSBL'  R5sx\��zRIENTTOp!C�oP�a.A�[ UT_SIM_ED��b�b[ V_ ?LCT z?�*�+^�)�_PEX9E�,&RAT8 jv�2u�p0"� UP ){.�PS0��/�/X�/�/�)�$O�2 ��m)deX)dh}��X d�� ?-???Q?c?u?�?�? �?�?�?�?�?OO)O@;OMO_OqO�O�H2
? �O�O�O�O�O__1_C_U_%�<�O_�_�_ �_�_�_�_�_o!o3o�Eo�O� �Ov 1r(���(���07�, ��lp�` @D� M �a?��c�a?m��a%�D�c�a���l�;�	l�b	 ��xJ��`�o�u��` �< �	p�� �r��H(���H3k7HSM5�G�22G��ޏGp
��������Yk|��CR�>���qȋs�a����o*  ���4�p�p��pT����B_����j�%��t�q� )�/��aD�������6  ���P�� Q� �� |��������	'� �� ͂I� �  ��i�=�������a�	���I  �n @)��mC�D��m��[��N���  '� ��~q�p�C�C�@�s�pC����ҟ 5�
�T�=x@#�7~9�$^�n�B�I�A��Q���� 0�q��bz 比������ȯ�����( �� -݂*�΁6����Am� �0rx���m�lp �?�ff U ܫN�`����Dn�8m྿̺>�'  P�aզ(m�������� q�c�d#?���m�xA�n�<�
6b<߈;�܍�<�ê<� <�&1j�m�A0��c���n��?fff?0�?&�����@�.�?J<?�`��l� ����dѩ�e�ϟg� ���d��Q�<�u�`ߙ� �߽ߨ��������)�  �M�8�q���
��j����f�E�� E�~0�G+� F�� ����� �F�1�j�U�P��y�[bB��A�� |����t�z���3 ��T��{�����<�t��h��u�w�>��*�N09K���A��Z��_�Cq�mc��?��//D///T)����pٞ�a�`CHT/A
$� !�!�@Iܝ�'�3�A�A�AR1�AO�^?�$��?�����±
�=ç>�����3�W
=�#�\>��+e�� �������{����<���.(�B��u��=B�0�������	3�\*H�F�G����G��H��U`E���C��+�Y-I#��I��HD��F��E��R�C�j=�>
�I��@H�!�H�( E<YD0X/�?O�?/O OSO>OwObO�O�O�O �O�O�O�O__=_(_ a_s_^_�_�_�_�_�_ �_o�_ o9o$o]oHo �olo�o�o�o�o�o�o �o#G2kVh �������� 1�C�.�g�R���v��� ��ӏ��Џ	��-�� Q�<�u�`�������ϟ ���ޟ��;�&�8�tq�\�(�����,�����]��������p!3�8�x��ӯp!4Mgs����IB+�+��a���{�E� E���s�����Ϳ���%Pe�P��(��{�4��I�[�իR�}Ϗ��ϳ�������  ���˿I�7�m� [ߑ��H� ߿�����������"�84�F�X�  m�������������2 �F�$�Gb���ϲ����!C���@�s����� �F� Dz/��� F�P D�!����������,>P�?��W�@@W
}����������
 W���� &8J\n�����*� ���˨��1��$PAR�AM_MENU �?q���  DE�FPULSE��	WAITTMO{UT+RCV/� SHELL�_WRK.$CU�R_STYL �G,OPT]�]/P�TBr/l"CB/R_DECSN ��, �/�/�/
???)?R? M?_?q?�?�?�?�?�?��USE_PRO/G %�%�?#O.�3CCR ���6G_HOST �!�!;DxO0JT �BO�C[OmA�C�O>/K_TIME"�B��  �GDE�BUG�@��3GI�NP_FLMSK��O(YT��9_*UPG�AUP \��g[CyH6_'XTYPE����?�?�_oo #o5o^oYoko}o�o�o �o�o�o�o�o61 CU~y���� ���	��-�V�Q��c�u���*UWORD� ?	{]	R}S��	PNSW��V$ڂJO�!���TE�@�VTRACECTL 1|q�� ��/ ���4���DT Q}q��c�(�D � � L� p�M�t�� v�O� �7���� @��� ������p�t�Qt�V�v�t�t���v�t���v�� v�t�t��v�N�v�!t�"t�#t�'�v�U%t�&t�'t�(t�E)t�*t�@�v�,t�U-t�.t�/t�0t�U1t�2t�3t�4t�U5t�6t�7t�8t�U9t�:t�;t�<t�=t�>t�?t�n v�@]�v�� v�� v�Dt�DZ v�Ft�Pv�Ht�It�Jt��Pv�s��������Q������ဨ�� ��U��V��W���X��Y��Z��[���\��]��^��_���`��a��b��c���d��e��f��g���h��i��j��k���l��m��n��o���p��q��r��s���t��u��v��wʜ�x��y���� ���&�֘�;Ҙ� #Ҙ�KҘ��P��� ��T� ������	��U
��������E�����@��������۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y���l�Е�� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_Е ���_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� ��_@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/�L/^/h!�$PGT�RACELEN � g!  ���f �|&_�UP ~��e��!� �!� �|!_CFG F�%�#f!�!��$�� �/�/;�"DEF�SPD ��,l1�� �| IN� �TRL ��-�f 8�%G1PE_C�ONFI� ��%O��!�$<WLID�#��-�4?GRP 1��7�!��g!A ����&fff!A+3�3D�� D]� CÀ A@6
B1�f d�$I&I�1~�0� 	 ?8�"�+@O ´yC[ODKB|@�A�OmOO�O��O�Of!>�T?��
5�O4_F^0_ �=��=#�
 K_�_G_�_�_�_�_�_�c_�_&o�_6o\oGo G Dz�c�of 
qo �oao�o�o�o�o0 T?xcu������IK
V7�.10beta1��$  A��E/�ӻ�A �f ,�?!G�C�>���+���0T�{��+�BQ�c��A\i�T�D;�{�p
�"�B������Ə�؏�T�O'O�2 �8��\�G���k��� ����ڟş���"�� F�1�V�|�g�����į ���ӯ���	�B�-� f��ov���K������� �����>�)�b�M� rϘσϼϧ������=�F@ ��'� ۫%Wك�W߉ߛߑ6 ���������%�� I�4�m�X��|��� ���������3��W� B�{���x��������� ����S~�w �8����� �+O:s^� �����
�<�// R�d�v�l/~/�ߥ/�� ������/�#?5? ? Y?D?}?h?�?�?�?�? �?�?�?O
OCO.OgO RO�O�O�O�O�O�O�O 	_�O-_?_jc_u_$_ �_�_�_�_�_�_�_o o;o&o_oJo�ono�o �o��(/�ob/P/ &Xj�/��/�/�/ �/��o��3�E�0� i�T���x�����Տ�� ҏ���/��S�>�w� b�������џ������ �+�V_O�a����p� ����ͯ���ܯ�'� �K�6�o�Z����o�o �o޿*<nD� rk�}Ϩ����� �������
�C�U�@� y�dߝ߈��߬����� ����?�*�c�N�� r���������0� ��;���_�q�\����� ������������7 "[F����ο� ���(�0^�W i�Ϧϸ�v�r� �/�///S/e/P/ �/t/�/�/�/�/�/�/ �/+??O?:?s?^?�? �?�?�?�?�?�O'O �?KO6OoO�OlO�O�O �O�O�O�O_�O_G_ 2_k_����_�_� 
ooJCoUo� ���oL_�o�o�o�o �o?*cu` �������� �;�&�_�J���n��� ��ˏݏO��7� "�[�F����|����� ٟğ���!���W� �_�_�_�����_�_ o����6b�$PLI�D_KNOW_M�  bd��j�#�SV �3e=�:e��z�����7�¿�������j�vmC�M_?GRP 1�P��`Ud�bd@I�߶
B�_�
�_����� t��@ǘϾ�^����� �Ϫ�
�����F��d� (�Zߠ�^����ߔ߶� ���*��� �f�$�L� ��Z�|���������X,�>�#�MR'É.�1Tg��� 㢞� ���������������� ��Q+%7��� �������M '!3��������Y�ST'�1 �1�3e3 �i�0:o A >/g�</ N/`/r/�/�/�/�/�/ �/�/?C?&?8?y?\? n?�?�?�?�?�?	O'�2(.:/j��<=O.3'O9OKO]O!#A4vO�O�O�O!#5�O�O�O�O!#6_&_8_J_!#7c_u_�_�_!#�8�_�_�_�_!#MA/D  wd3#x`�$PARNUM � ++�5o"S+CHOj ]e
�gpa8�i=��eUPDpo�e��t"_CMPa_$�R`ؠ`';�~)tER_CHK7u���;�Or4F{RqS|�2�#�_MOQ`��u_�be_RES_G' �+-O� ��H�;�l�_����� ��Ə���ݏ����w&@�|�5��uu@ R�q�v��s�@������ �sPП����sbP� .�3��s�PN�m�r��s� `�������rV 1�P���b@cX���p�$@cW��(��(�@@cV��4���rTHR_ICNR|�Taud<�oMASSI� Z]��MNH�{�MON_�QUEUE ��.�bvg��g�bdN�.pUrqN��`{ΰE�NDб��EXE����`BE��ڿ˳OPTIO׷�{ΰ�PROGRAM %��%Ͱ믖o~̲TASK_IQd�@�OCFG �𮿄o����DATA�e���@�2 �N�`�r߄ߒ�<ߵ� �����ߖ��!�3�E�W�
�INFOe�"ݘ��������� ����)�;�M�_�q� ��������������hn�z�"� !����OpDIT ����s�WERFL���#RGADJ7 �b
A��0��?��P��IOR�ITY��av��M�PDSPX��U�����OG$ _�TG� K���ETO�E��1�b (/!AFD�E�p�~�!tcp�>�!ud��?!icm��F�XY_���b=���)� *J/\/` ���G/�/k%w/ �/�/�/�/�/?�/2? ?V?h?O?�?s?�?�?=*�PORT3�Rc����u�_C?ARTREP�b>k@SKSTA���z�SSAV���b
	�2500H86A3(�ς5D1�b`@�����s�Ox�O�G	PURGE��B�	�yWF�@DO��$�evW�T�a�:�WRUP_DEL�AY �bTRO_HOT{��%o��_TR_NORM�AL{�}_�_�VSE�MI�_�_oCaQS�KIP1��u�Cx 	bO\o\@Jo �o�o�ojh�u�o�g�o �o	�o?-Ou ��_����� ��;�)�_�q���I� ������ݏ��Ǐ%� �I�[�m�3�}������ǟٟ�ͥ�$RB�TIFR�RCV�TM.+D�	�DkCR1c�8l�qi�C ��>�� �>�k��o �U	��I�i���nro¯��<�
6b<߈;�܍�>u.�?!<�&ǯ ���)�ŰHB�T�f� x���������ҿ��� ���>�)�b�Mφ� qσϼϟ�����5�� (�:�L�^�p߂ߔߦ� �������������6� !�Z�E�~��s���� 	������ �2�D�V� h�z������������� ��
��.RdG ������� *<N`r�o �����/�&/ 	//\/��/�/�/�/ �/�/�/�/?"?4?F? X?C/|?g?�?�?�?�? �?�?�?O0Os/TOfO xO�O�O�O�O�O�O�O __,_OP_;_t___ �_�_�_�_�_�_oGO (o:oLo^opo�o�o�o �o�o�o�o�_�_$ H3lW���� �o�� �2�D�V� h�z�������ΈB��GN_ATC 1��O� AT&FV0E0΋�ATDP/6�/9/2/9��ATAΎ,�AT%G1%B9�60�+++�3�,.�Hc�,B�I�O_TYPE  �����ЏRE�FPOS1 1�>�� x��������?�P���� 6�������V�߯z��� �9�Ǜ2 1�����$��� �ƿ<D�ё3 1�^�p������:�%�^�ܿS4 1����Q��������q�S5 1� �ϚϬ���d�O߈��S6 1��/�A��{�������S7 1���������y�|��0�S8 1�G�Y�k��#��G���SMASK 1����  
����e�XN	O��;�A�����͑?MOTE  ��ʔ���_CFG ����<���̒PL_R�ANG���q��PO�WER ���^ ��SM_DRY�PRG %��%���dTART ��V�
UME_�PROs� ʔ_�EXEC_ENB�  =���GSP�D� #��4TD�B>PRM_PMKT_m�TQ �����OBOT_NAM/E ���׉�OB_ORD_N_UM ?V���H863 � �t ��e!\<�  #� 	r*!@��"D|<���PC_TIMEOUT6{ x��S232
�1�� L�TEACH PE�NDAN_ ����e����Mai�ntenance Cons�r���*�"�/�KCL/)C� :���/?� No Us�ee��/U?�v#NPqO218����t!CH_L� ����7�	�1�;MAVAIL�a#��������SPACE�1 2�ٜ ��?%dH�9�eF%��<��L8�? H �9�O�?�O�O_�O (_#WTOfOxO�O8_�O �O�_�_�__o i� �4mT_f_x_�_�_�_ �_�o�o�oo .�5;A2@NROdovo �o6�o�o����4��I�N{3]o� ��S������ޏ 0�Q�8�f�N{4z��� ����p����8�@��M�n�U���N{5�� ����͟ߟ���%�4��U��j���r���N{6 ��Ưد����� �B� Q�r�5χϨϏϽ�N{7ѿ�������=� _�nߏ�Rߤ��߬���N{8�� ��$�6��� Z�|ߋ��o���������N{G ���� ���$
�� C�e#p��������� ����:hL���2��+��^�!dt Y�k�� ������� 8oR~q�� ����//=/ 7Ikm�/���/ �/�/??+?=?3/]?pW/i/�/�= `�� @NP�5<�?�/�) A�5�?1OCOI? #J$OVO�O�O�O~O�O �O_�O�O�O_^_ _ 2_D_v_�_�_�_�_�_ o$o�_�_
o<o~o@o�N<
O�oN{_MO�DE  +��iS �+��ox?v:A_��?'y�z	���o�CWORK_{AD�mvτq�/R  +������p_INTVA�L�`@�zR_O�PTION1� �u��VAT_G�RP 2�+�]�(���L��ԏ揥�
�� .�@���d�v���O�o ���dX�ß����ϟ 1�C�U�g�)������� ��ӯ�{�	��-�� �c�u���I�����Ͽ ��ϛ��;�M�_� !σϕϧϹ�{����� ��%�7���[�m�� Aߏߵ����ߛ���� !�3�E�W���{��� ��s����������/� A�S�e�w�������� ������+��O as���?�� ��'9K[�����e�$SC?AN_TIM�a���\��R �(�30(�L8z�_�p�p	
WtZ��2#Nq!»#Y�:.(/1��#M"2{$!!d��(~!�!�r #]) �0��/�/�/�r�)�/�  P5�0�2  8�?U?g?>1D��j?�?�? �?�?�?�?�?O#O5OpGO?Nq�%ROЌO�O[N![q;��o�t�Nqp]M�t��Di�t|!c{  � lM" Nq�A!
%�1_C_U_ g_y_�_�_�_�_�_�_ �_	oo-o?oQocouo �o�o�o�gS�o�o�o '9K]o� �������� #�5�G�Y��o�o�K�� ����Џ����*� <�N�`�r����������̟ޟ����1�  0�B|�_g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ�p���)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑ��ϐ����� ����0�B�T�f�x� ���������������,�>�P�J�V�   �1�������������� ��1CUgy �������	 �y3"HZ l~��������C&5/</+&��r! 5/q-	�1234567}8R���L{0�@�/�/�/�/�/?3,?>?P?b? t?�?�?�?�?�?�?' OO(O:OLO^OpO�O �O�O�O�O�?�O __ $_6_H_Z_l_~_�_�_ �_�O�_�_�_o o2o DoVohozo�o�_�o�o �o�o�o
.@R dv�o����� ���*�<�N�`�� ��������̏ޏ��� �&�8�g�\�n����� ����ȟڟ����"�+&s�C�U�:�Z���������Cz  �Bp   ����2/$@��$SC�R_GRP 1��(�e@(�l��� @� Z! �U!m�	 #�-�=�6�n�p� l�S�y(J�w�e�����7�3%Dʰ֠�o��ป���M-10iA 890�%90� Ɓ ?M61C �#�-�I���#�
\�l� ,�O'|�Z!�S�;�o�}�	n�����������X �,���Y" N�a����ߖ�i�@�.!�`/��m�����"��B�Š�J�H�a�H�9A֠p�  @. ��Dl��?���D�HŠ����H�F@ F�`�������;� &�K�q�\�������<퀈����������B���YD}h� ������
 CҾ?4#��0/v/�%���
������3�V�j�@���/7 B�*'���P���EL_DEFAULT  CԿ����X!MIPOWERFL  P�p%W"�} WFDOe& �p%��ERVENT? 1���I�n#�=�L!DUM�_EIP��(�j�!AF_INExd ?�!FT�/�7>�/[?!K߀? ��J?�?!RP?C_MAIN�?�8q��?�?�3VIS�?�9��??O!TP&2@PU6O�)d.O�O�!
PMON_POROXY�O�&ezO��ORB�O�-f�O#_!RDM_SR�r�*g_o_!RL(d�_�$h^_�_!
�0�M�O�,i�_o!?RLSYNCo.i�8�_So!ROS�/zl�4Bo�on? �o2S�o�o�o�o5 �oY }D�hz �����1�C�
��g�.���R����'ICE_KL ?%�+� (%SVCPRG1������D��3$�)��4L�DQ��5t�y��6�����7ğɟ�=��/�9��脆_A� ��i������>� ���f��끎�	�� ��1��ޟY����� �.����W�ѿ�� �����!��ϯI�� ��q������G��� �o���������� 9�;�翹�˂�ҏ� ����á������� � 9�$�]�H���~�� ����������#��5� Y�D�}�h��������� ������
C.g R�v����� 	�-QcN� r������/�)//M/��_DEV� �)�M{C:U(��]g$OUTYB`!x&c(?REC 1���` �  `  	� ` ` ` @` �!�!U+�#��U/�.�$1�"?`!�` 8:
 ��P�b6 �s�'�  ��  '� �  =0f���"�#�!U� ` /` �` ���=y �y �y ������` B� D��?O�%��|0��<S7  ��H� �0�_��? O�U` �4)` ��?S��`!y ��0�` �k� NPO�OOc�ʀ;[0�0�1o�  �� i�O U!� � �04,` -�xO��y ��!�D�n� M�O]_�Oc��O�@�F��O
__�._@_R_d_If�6Wr _�H�i@�4��x�C�@��_�!�r` �` C` �P�#�_�fy �y �
y �y �<1To�oo�h$0k �  �� �1   �
i@=�o ;@�2�0� �  K`$|o�dJy �y �y Dq��!X a�oh[�l�0|k`�bR  Ȣ QlP
5�2` �` ��(�c�4��D�p�!��t~�j�0km� ��3��`�  #"�j2;*� ` L` �� wOW���y �y ��q�y ��QX���ta��<Đ?g���?�?��?�?��ď"F �;�T�f�4���'��+�` =� �� ��
j` Q� ,�����U�H��` U� F�� �x�02y0 � �T�B� x�f�������ү��� ���,��P�>�t��� h�����ο��޿�� (�
�8�^�Lς�pϦ� �����Ͼ� ���$�� 4�Z�H�~�`�rߴߢ� �������� �2��V� D�f�h�z������� ��
���.��R�@�b� ��j����������� ��*<`N�r�����%V 1͸�, P 8� :����*��o 
GxS�Jc(TYPE�/�e"HELL_CF!G���&� ��"�>� %RS�p� ��//?/*/c/N/ �/r/�/�/�/�/�/? �/)?8;�p:>����` %K?y?�?F=J1�J1�p gA�=�1�p)��a22!�d�?�?��HK 1�� �a�?AO<ONO`O�O�O �O�O�O�O�O�O__�&_8_a_\_n_�_|OMM ���_FTOV_ENO��nwOW_RE�G_UI�__IMWAIT�Rq�6k�OUTf iT�IMe��ZoV�Aw�1o#a_UNI�T�S�fwMON_�ALIAS ?e~�Y ( he �o�o0��o] o��>���� ��#�5�G�Y�k�� ������ŏ׏����� �1�܏B�g�y����� H���ӟ���	���-� ?�Q�c�u� ������� ϯᯌ���)�;�� _�q�������R�˿ݿ ��Ͼ�7�I�[�m� �*ϣϵ����τ��� �!�3�E���i�{ߍ� �߱�\��������� ��A�S�e�w��4�� ���������+�=� O���s���������f� ����'��K] o�,����� �#5GY} ����p��/ /1/�U/g/y/�/6/ �/�/�/�/�/�/?-? ??Q?c??�?�?�?�? �?z?�?OO)O�?:O _OqO�O�O@O�O�O�O �O_�O%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3o�_Woio{o�o �oJo�o�o�o�o�c��$SMON_D�EFPRO ����4q� *SYS�TEM* . �"vRECALL �?}4y ( ��}7xcopy �fra:\*.*� virt:\t�mpback~q=�>desktop�-b25t4o0:15916 �q����y}
xy�zrate 61 ��4�F�X��u� �w�8360 @�'���ʏ܏o�1}�@����2�D�V��w6ur�md:program_1.tp�emp\���+��� Οa�s�����:�L� ^��{��#���Ưد<���:544���� 6�H�Z�����#��� ƿؿk�}�������<� N��󯅿��)Ϻ������ }:uts:o�rderfil.dat�~Ϧ�/�A�4S�f�1��b:��@��&߷������r5tu�}��Ǫ�;�M�_�}6t�� +���� a���ߎߩ�:�L�^� q����'��������� ���%�6HZm��� ��������� !�2DVi�{��� ��������./ @/R/ew/�-/�/ �/���/�/<?N? �/s?�)?�?�?�? ��/�?'/8OJO\Oo/  OO�/�O�O�Om�O@�O�O4_F_X_�E!t��432 _(_�_ �_�_pY|��_�_1oCo�Uo�H7���o2  ,o�o�o�_t_o�o ;M_�_�(� ��po�o~�7�I� [��o��$���Ǐُ l~�����3�E�W�� �� ���ß՟�z�@���/�A�S��*;�/�?�������ӯ�*2 t?�����8�J�\�� ��$SNPX_A�SG 1������� �P 0 '%�R[1]@1.Y1`���?��#%�� ֿ����ݿ�0��:� f�Iϊ�m���ϣ��� ��������P�3�Z� ��iߪߍߟ������� ���:��/�p�S�z� ������� ���
� 6��Z�=�O���s��� ���������� * V9z]o��� ��
��@#J vY�}���� /�*///`/C/j/ �/y/�/�/�/�/�/�/ &?	?J?-???�?c?�? �?�?�?�?�?O�?O FO)OjOMO_O�O�O�O �O�O�O�O�O0__:_ f_I_�_m__�_�_�_ �_�_o�_oPo3oZo �oio�o�o�o�o�o�o �o:/pSz ����� ��
� 6��Z�=�O���s��� Ə���͏ߏ ��*� V�9�z�]�o������� �ɟ
����@�#�J��v�Y�r�PARAM� ���� ��	�z�P���j�OFT_K�B_CFG  �����ѤPIN_S_IM  �Ʀ��)�;�ɠr�RVQSTP_DSB ��Ƣw�����SR ���� & 胿����ΦTOP�_ON_ERR � ����PT�N ���AݲRINGo_PRM� ���VDT_GRP �1����  	 ʧ��\�nπϒϤ϶� ��������%�"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�w�t��� ������������ =:L^p��� ��� $6 HZl~���� ���/ /2/D/V/ h/�/�/�/�/�/�/�/ �/
??.?U?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo mojo|o�o�o�o�o�o��o�o30ѣVP�RG_COUNT�����^rEN�B)�YuM�s㤐_�UPD 1��8  
G���� �'�"�4�F�o�j�|� ������ď֏����� �G�B�T�f������� ��ןҟ�����,� >�g�b�t��������� ί�����?�:�L� ^���������Ͽʿܿ ���$�6�_�Z�l� ~ϧϢϴ�������VuYSDEBUGhp��p���d�y�SP�_PASShuB�?.�LOG �V�u�s������  ��q��
�MC:\Z�
�[�_MPC`��u�����q���� �q��SA/V �c��ԛҶ����SV�T�EM_TIME �1��{ (�p��t���s�N|T1S�VGUNS�piu'��u���ASK_?OPTIONhp�u��q�q��BCCF�G ��{I� 8B��5�`5�;z C�l�W�i��������� ������2D/h S�w����� 
�.R=va�������� /��B/-/f/Q/�/ �/�� �/�/�/�/ �/ ??D?2?T?V?h? �?�?�?�?�?�?
O�? O@O.OdORO�OvO�O �O�O�O�O_�H�_ ,_J_\_n_�O�_�_�_ �_�_�_�_o�_4o"o XoFo|ojo�o�o�o�o �o�o�oB0R xf������ ���>�,�b�_z� ������ΏL����� (��L�^�p�>����� ����ܟʟ�� �6� $�Z�H�~�l������� دƯ��� ��D�2� T�V�h�����¿x�ڿ �
��.Ϭ�R�@�b� ��vϬϾ��Ϟ����� ��<�*�L�N�`ߖ� �ߺߨ��������� 8�&�\�J��n��� ���������"�ؿ:� L�j�|���������� ����0��TB xf������ �>,bPr ������/� //(/^/L/�/8��/ �/�/�/�/l/? ?"? H?6?l?~?�?^?�?�? �?�?�?�?OO OVO DOzOhO�O�O�O�O�O �O�O_
_@_._d_R_ t_v_�_�_�_�_�/�_ o*o<oNo�_ro`o�o �o�o�o�o�o�o 8&\Jln�� �����"��2� X�F�|�j�����ď�� ԏ֏���B��_Z� l�������,�ҟ�������,��J��$T�BCSG_GRP� 2����  �J� 
? ?�  u��� q�����ϯ��˯���)�;�N�U��\�d�, �j�?J�	� HC��8�>󙚆�9�CL  �B�m�����z�ݸβ\)��Y g A���B�;�F�Bl�=�,�ɐ�|Z�,��  D	�{�F�`�j�Cs��ό�$�ϰ̖���@J�� +�>�Q��.�|ߙ�dߠv��������؈J�	V3.00m��	m61c��	�*,�$�I�;�D�>ə��J�(��� �r�D�s�  #�����D���N�JC�FG ���f� i������r������� 7�E��E�k�V���z� ��������������1 U@yd��� ����?* cN`����� �m����/"/�U/ @/e/�/v/�/�/�/�/ �/	??-?�/Q?<?u? `?�?�?J�6��?��? �?�?*OONO<OrO`O �O�O�O�O�O�O�O_ _8_&_H_J_\_�_�_ �_�_�_�_�_�_o4o "oXoFo|o�o���o�o bo�o�o�oB0 fTv���~� ����>�P�b�t� .���������̏Ώ�� ��:�(�^�L���p� ������ܟʟ ��$� �4�6�H�~�l����� Ư���د�� ��o8� J�\����z������� �Կ
���.�@�R�d� "ψ�vϬϚϼ����� ����<�*�`�N߄� rߨߖ߸ߺ������ &��J�8�n�\�~�� ������������ � "�4�j�X���|����� n���������0T Bxf����� ��,P>t ���d���� /(//L/:/p/^/�/ �/�/�/�/�/�/? ? 6?$?Z?H?j?�?~?�? �?�?�?�?�?OO O VO��nO�O�O<O�O�O �O�O�O_
_@_._d_ v_�_�_X_�_�_�_�_ �_o*o<o�_oro`o �o�o�o�o�o�o�o 8&\J�n� ������"�� F�4�V�|�j�����ď ������O�$��O�� f�T���x�������� ҟ��,����b�P� ��t�����ί௚�� ���(�^�L���p� ����ʿ��ڿ ��$� �H�6�l�Z�|�~ϐ� �ϴ��������2� � B�h�Vߌ��8����� rߠ�����.��R�@� v�d��������� �����N�`�r��� >�������������  J8n\�� ������4 "XFhj|�� ����/0/��H/ Z/l//�/�/�/�/�/ �/�/??>?P?b?t?�2?�?�?�?�?�?�> s @
C 
F�O
B�$TBJO�P_GRP 2���5� � ?�
G6B=C��DL��0�_xJ�@�
D�@ �< ���@�
D @�@UB	 �C��} �Fb  C�VG<UAUA>����E�E��I>��@�A�33�=�CL�@f�ff?�@?�ff�B�@Q�E-_8W�N���O>�nR\�)�O�@�U���;���hCY�@� � @�@UAB�  �A�$_�_�S�UC�  D�A�LwP�R�O�z_�Sb��
:���Bl�P���P�D�Q�_So
AA�ə�A�hcZQD9Xg�F�=q�e
o��@�p��b�Q�;�AȰ@�o��@L�CD	x`��`�o�ojo|o>B��\u�oh�Qts>�a@33@QV@C��@�`ew�o�>��D�u*�@�x p�qP<{�Nr�@@�PZv_p��� �&�:�$�2�`���l� &���ʏ����!��� ��@�Z�D�R�����DT�
Fґ�E	V�3.00�Cm61c�D*���DA�
�� Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I&�CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;'`�;Q���8�`�F�O���
F���Q��K�2DESTPARS  �8�O@3CHRe�ABL/E 1�DK.�
C�P�%� ~ �P�BP�P�	GAP�	P�E
P�P���
AP��P�P�|�RD	I��NA����¿Կ���`�Oh�z˄ϖϐ�Ϻ��΀�Sf�LC  *ʍߟ߱��������� ��/�A�S�e�w�� ��������)Me�i� ��$���1�C�����%�7�IȀ�
�NUoM  �5NA�@@ ��[���_CFG ������A@6@IMEBF_TTk���LCx��5VERY�6�K�5R 1�DK
 �8�
B@� �0/�  ���� ��� 2DV hz�����/ �
/S/./@/V/d/v/Ru_��b@L
6@MI_CHANA� L �#DBGL�VPCL5A� E�THERAD ?U�550�M��/��/N?0F� ROUT6_ !DJ!�4�?~q<SNMASK*8|LC;1255.�5���?�?2DOOLO_FS_DIk��%�9ORQCTRL� �mK���hM8 WO�O�O�O�O�O�O�O 
__._@_�|ON_`_��_a�PE_DET�AI8-JPON_�SVOFF#O�SP_MON ��J�2�YSTRTC_HK �DNg?��RVTCOMPA�T�X53�T�PFPR�OG %DJ%	>qaRAM_17o�\�APLAYl��Z_�INST_M�0 2�l�W�dUS_Wo�ibLCK�l�kQUICKME� #iboSCRE@p-:tps�ib�a[p`y�"qp_uy��Ti�9SR_GRP �1�DI ���0��z���5�#�Y�G��2 ���� S��o����܏ǅ��� �)��M�;�q�_��� ����˟���ݟ���7�%�G�m�	1234567堃����b�XZu1��{
 ��}ipnl/�ՠgen.htm������*�<�R��Panel s/etup@�}6o��`������ȿڿ o� e��$�6�H�Z�l�� ��ϴ���������� �ϗ�D�V�h�zߌߞ� �C�9�����
��.� @��d��߈���� ����Y�k��*�<�N� `�r����������� ����8��\n�����-�nUA�LRM�`G ?DK
  �	 L?pc��� ����//6/��SEV  ��h&�ECFG ���]�&��A�! �  Bȣd
  7/�c-5�/�/�/?? %?7?I?[?m??�7t!�r��[ �3ȏ�?�B'Imf?wk�P(% */O`
OCO.OgORO �OvO�O�O�O�O�O	_0�O-_�<�d �=�?�;_I_?pHIST� 1��Y  �(�  ��(/�SOFTPART�/GENLINK�?current�=menupag?e,153,�o�_x�_oo �� �_�]936�_lo~o�o �o1b�o�o�o�o %�oI[m�� 2�����!�� E�W�i�{�������@� Տ�����/���S�@e�w����������L� �QL������1�C� F�g�y���������P� ���	��-�?�ί� u���������Ͽ^�� ��)�;�M�ܿqσ� �ϧϹ���Z�l��� %�7�I�[���ߑߣ� ������ğ֟�!�3� E�W�i�lߍ����� ����v���/�A�S� e�w������������ ����+=Oas ������ �'9K]o� ���������� 5/G/Y/k/}/�/��/ �/�/�/�/?�/1?C? U?g?y?�?�?,?�?�? �?�?	OO�??OQOcO uO�O�O(O�O�O�O�O __)_�OM___q_�_ �_�_6_�_�_�_oo %o/"/[omoo�o�o �o�_�o�o�o!3 �o�oi{���� R����/�A�� e�w���������N�`� ����+�=�O�ޏs� ��������͟\�����'�9�K�6o��$�UI_PANED�ATA 1�������  	�}]�����0ȯگ��� ) �$� ᔒ�O�a�s������� �Ϳ�����'�� K�2�oρ�hϥό���p�������� Ha$�7�<�N�`�r߄� ���Ϻ�-������� &�8�J��n�U��y� ����������"�	��F�-�j�|�c���� ����������+ =��a�߅��� ��F�9  ]oV�z��� ��/�5/G/���� }/�/�/�/�/�/*/�/ n?1?C?U?g?y?�? �/�?�?�?�?�?	O�? -OOQOcOJO�OnO�O �O�O�OT/f/_)_;_ M___q_�O�_�_?�_ �_�_oo%o�_Io0o moofo�o�o�o�o�o �o�o!3W>{ �O _�_����� �pA��_e�w����� ����&����܏� � =�O�6�s�Z���~��� ͟���؟�'��� ]�o���������
�ۯ N����#�5�G�Y�k� ү��v�����׿�п ���1�C�*�g�Nϋ� �τ���4�F���	�� -�?�Qߤ�u߇����� ���������l�)�� M�_�F��j���� ��������7��[�����}�l�������������)��$�� Pbt���� ����(L3 p�i������ /(�����$UI�_PANELIN�K 1����  � � ��}1234?567890Y/k/ }/�/�/�/�$��W/�/ �/??+?=?�/a?s?@�?�?�?�?S9S *4�=��U   �?O (O:OLO^O�?\1O�O �O�O�O�O�O�O_(_ :_L_^_p__~_�_�_ �_�_�_�_�_$o6oHo Zolo~oo�o�o�o�o �o�o�o
2DVh z$�����
�E0,/A�M�/� p�S�������ʏ܏��  ��$�6��Z�l�O� ���<�?�����T!� ��1�C�U�g�Z3�� ������ǯٯ�z�� !�3�E�W�i��<���� ����C��ÿտ��� �Ϥs5�G�Y�k�}� �ϡ�0���������� ߮�C�U�g�yߋߝ� ,���������	��-� ��Q�c�u����:� ��������)���M� _�q���������(��� ��~���7I,m b������ �3ƞ����՟w� �������/�� ,/>/P/b/t/�//�/ �/�/�/�/??���� ��^?p?�?�?�?�??� �?�? OO$O6OHO�? lO~O�O�O�O�OUO�O �O_ _2_D_�Oh_z_ �_�_�_�_�_c_�_
o o.o@oRo�_vo�o�o �o�o�o_o�o* <N`����� ������8�J� -�n���c�����ȏڏ I��m"��F�X�j� |��������/֟��� ��0���T�f�x��� ����?/?A?�o�� ,�>�P�b��o������ ��ο�o���(�:� L�^�p����Ϧϸ��� ����}��$�6�H�Z� l��ϐߢߴ������� �ߋ� �2�D�V�h�z� 	�����������g �.���R�d�G���k� �������������� <N1r��� �;��&8J =�n������ i�/"/4/F/X/ǯ ٯ믠/�/�/�/�/�/ ?�/0?B?T?f?x?�? ?�?�?�?�?�?O�? ,O>OPObOtO�O�O'O �O�O�O�O__�O:_ L_^_p_�_�_#_�_�_ �_�_ oo$o�_HoZo lo~o�o�o��o�og �o�o 2VhK �o���������o�/�/�u��$�UI_POSTY�PE  �%� 	e������QUICKMEN�  ��d�����R�ESTORE 1�ݏ%  ���,�>�b�m]���������Ο q����(�:�ݟ^� p�������Q���ůׯ I��$�6�H�Z���~� ������ƿؿ{����  �2�D��Q�c�u�� ���������ϛ��.� @�R�d�߈ߚ߬߾� ��{υ����s�%�N� `�r���9������ �����&�8�J�\�n� �{������������ "��FXj|� �C������oSCREր?ۍu1sc'�Wu2G3G4GU5G6G7G8G��USER).@�T(IksQ�4��5�6�7�8����NDO_CFoG ޖ�  &�� ��PDATE� ��N�one V��SE�UFRAME  ���&!RTO?L_ABRT1/���H#ENBR/C(GR�P 1���Cz  A��#�!�@�/�/�/�/�/ 6
?�?A*ՀUr(A!a+MSK  u%}1a+MN.!%[�~2%���?��VISCAN�D_MAXs5I��](�0FAIL_�IMGs0`���#�}(�0IMREGN�UMs7
�;BSI�Zs3&���,~CONTMOUQ �u4��PE��c�� �@��"�FR:\�? �� MC:\�RC\LOG�FB@� !�?�O�A�O�_�z M�CV�O�CUD1&*VEX3[�`�qF��"ᖉ�`(��=7��͍_��Z�_ �_�_�_�_�_�_oo�,o>oPoboto�o�;P/O64_9C�B ��gn6�eK LIA��j�h�aV��lfy@�g�o� =	�hwSZV�n����g�WAI�o�4STAOT �+�@�O���z$���5J!�2DWP  ��P G)����a��;@'��2_JMPE�RR 1㖋
 � ��2345678901|������� ď��ɏ����B��5�f�Y�k����<N0M�LOW{~�@�0�@_�TIYH�'�0M�PHASE  �%���3SHI�FTO21"x[
 <���?\��;�a� ��q���Я�����ݯ ��N�%�7���[�m� ������ɿ�ٿ�8�@�!�n�E����*	VSFT1�c�V�0M�� �5ԩq� � ��EAȯ  B8�����"� p�����ª��B F��ME$�u4���\�a{~&%��M�i�x[�p�30�$xpTDINEND]H^8t�Or0U?��[J���S�ߏ���s5����Gy�	��,��������ߍ�RELE� �s/q�XOjFt�_ACTIV��~8��
 A �;}�<����RD�`��C!YBOX �����v���p2��>�190.0.���83����25	4�����`��� �q�ro�bot�ę�  � pHa�upc���u��p���r���ZABC�#�-,u� �r �5X?Qcu �����/�0/�/)/f/�Z;D�q� ��