��  ҥ�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Z  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
FPCOU�PLED1 $�[PP_PROC�ES0 � �1���UREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$,NO/P�S_SPI_IN[DE��$DX��SCREEN_NAME �/SIGNj���&PK_FI� 	$THKY��PANE7  �	$DUMMY1U2� �3�4�~GRG_STR1� � $TI�T�$I��1�&�$�$�$5�&6&7&8&9'0''�%!'�T%5'1?'1I'1S'�1]'2h"�ASBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGW�~0�$	Y $DB\� � COMqW��MOJWH.
 �\�VE�1$F8 �A�$O��D��B�CTMP1_F�E2�G1_�3�B�2�H X_D�#� d $CA�RD_EXIST��$FSSB_�TYPitAHKBgD_S�B�1AGN �G� $SL?OT_NUMZIQOPREV��G ��1_EDIT1� � h1G=�H0S?@f%$EP<Y$OPc ��0LETE_O�KRUS�P_CRQ$�4�VAZ0/LACIwY1�Rp@Pk �1w@MENP$D�V�Q�P�ЩA��nQL*OUyR ,lA�0V1�AB0~ OL]eR�"2CAM_;1� x�f$AT�TR�MP0ANN��@�IMG_HE�IGHQ�cWID�TH�VTC�U��0F_ASPEC�Q$M@EXP�;�@AX�f�CF�T X $GIR� � S!1�@B`�NFLI�`t
U�IREs3�tGITSCH~C�`N.0S�d�_L�`�C�"�`E�Dkp;tL0J*DS��0>0�zra4 gq;G�0 � 
$WARNM'@f�+P�� �s�pNST� C�ORN��1FLT�R�uTRAT@0T��p  $AC�C�1
� ���OcRI	`!S<{RTq0�_S�B�qHGI.1 [ Tpu3I8�TYVD+P*
2 �`v@� 1R*HD�cJ* ���U2��3��4��5��U6��7��8��9�;CO�$ <� �#5x�s1v`O_M|�@�C t 0�Ev�NG��ABA� �c��YQ�������@������P��0����x�p��PyP�2� ����J��_R��BC�J���2�JVP�C�R��}@w��u�tP_�}0OF� 2  @�� RO_����aIyT8C��NOM_�0r�1åq3��T �#���@xP��J}EX�G�0�� .��p�
$TyF`��C$MD3���TO�3&@U=0�� ��H�2�C1{�E͡� vE�uF0�uF��0CPo@�a�� 	P$@`PU8�3�f)"��&)�AX 1rDU6�$;AI�3BUFV�@Ȳ�! |�pڶ�p[PI��PZ�EMY�Mf�̰i�FZ�SIMQS��/�ȩA-�����kw 	Tp{zM��P�B��FACTqbGPE�W6��Ҡ��v��M�Cc� �$}1JqB�p;�}1DECG����G��A-�b� ���0CHNS_EMP��$GO���+P!_��q3�p�@Pۤ��TC��{r��q0�s�� a�/�� �B���!	����JR!0��SEGF�R��Iv �aR�TrjpN%S+�PVF�����ʹY�K���a1�)B���( 'j�Av�u�ct��a D�.0���*�LQ��DчSIZC������T���O�����aRSINF�����jq��C��C����LW������x�CRCLuFCCC kpy�����N}���b�A�������d��D
wIC��C���r��+ 0P��z�2EV2�zUFH_��FpNt�/�>����rH�1Q��!  ��@ �Qx����U�kp�2 ݠ�a��s�+����R>T!x "�4��4u2��tAR���`CNW�$LG�p��B�1 �Pr�P�t�aA?@z��ϣ~0R�ӲME`�`8�oC�RAs3��AZ����pb�OFS�FC�b�`�`FMpp�� �0��ADIS+ �aV%��b�z��pE$�pRp�cV�S�P��a&+QMP5�`Y8C��IMe�pU��aUSw" $=�TIT�1��S�SG1��#�8��?DBPXWO! T=#��$SK��2��DBTmTRLS$l�Q0TQ��P`�P�D�q�1LAY_CAL�1�R^0o f7#PL)A�Q�D'a�7�3a�7��(3!S%�2?�PRj� 
p*0���S& =�6A$��$ �*ЅL�9'�?'�U�T(�O�A�PCS)�#ODENE��1*BO'Ӳ0RE�pB_+H �Ou�o&$L�C'$�3�R��K2�LVO�_9D~!U�ROSbrq��v�R����CRIGGER�FPA�S��6�ETURN�B�cM[R_}�TUbp���@EWM$���G1N=`���BLA��TU�ܡ($P�)$P s�*hP3a��1C�TΣ@DO>���D�A���FGO_A7WAY�BMO"�a��!*0CS_P,<aISt�� ��� �s�S#�Q����Rw�cV��Qw2�VW���'dNTV(��RV ;����~��mgŃ���Jt��<@��SAF�Eڥ�f_SV�bEOXCLUT��� 'ONL���cYfЀ��y�OTEuHI_�V} ��PPLY_|�q7�VRFY_b3����Rj L�_ -�h@0��_y�1� �o��QSG�  .�rŐ1PNQ5�� _q���;P��Vby|rsvANNUN<@�$�tKIDX�UR�c[P@� �y�qi �z�v)1�EF�PI<B/��c$F�r�$АOTQP��A $DUM�MY��&���&����*0t�U0 `  �HE�\���^r�c|YRr SUFFI����Pa0��P)�5�#�6#�)1MSW��U1 8��KEYI��4�TM�A��ځL3QՆINݱv����j P2 D��HOST�0!��������������EMp&����*0SBL� ;UL��3 Z����D�*0T�@S4 ϴ $���USAMPa༥.�������V I�@��$SUB����;@c����3��SAV�������������`�vP$�@EC!	0YN_Bn35 0��DI�tb�PO\�M��#$E��R_IB� �E�NC2_S�T6X��2������ �cG���0 S72��1���A����8  A��Ǜ��@PK�Dxk!uq��AVERҁ8�����DSP�ܢPC?���26�\������VALU�HE4 �M_�IP(�ܣ�OPP� 5�TH��ͫ��S` 4�.�	FB�6d��~�� 5��SC?q���ET��9ȂFULL_DU���qKP�ԝ�����OT�"T�P�NOAUTOS:��$YĪ�Z� �T��X�C�0h�CE2�6�1V�L� _;H *h�L� �����$P��wc �ě1�Ʃ1��C��Ƨ���Ʋ���7��8��9R��0����1��1��U1	�1�1#�10�U1=�1J�2X�2�˪��2��2	�2�2�#�20�2=�2J�3JX�3��3����3	�U3�3#�30�3=�53J�4X����;SE�2< <8�Z����I��e�$�}ōJpFE5P?PT=� ,f��a? ��P�?i��e�i�E�Pq���azT>F�$TP$!?$VARI���n�UP21p? 7���TD��s��p��t����	��BAC2@ T����$uP�*p��Þ0� IFIw�0�P� � )PB"�IqF0P�TAt� ;u�"�"pu STvt: �bt�@�Tl�6	sC2	>0 ���S���/bF���FORCEUP�sr��FLUS�pH�fNn����bD_�CM�PEv*I�N_t�e`�REM� F�a�a�0�(Te�KdN~�e�EFF�j�PIN�Ja�OVM�OV=A�TROV���DT	��DTMX ,A��P*��0M(�xR#�0�CL*_ ��u*�Pr�{_XЉ�_T�+X��PASaD% ��(װ�1�`�&_A@RQ�LIMIT_�4�� �M��CL�tˑR�IVW�*2EAR6�IOxPC�P��2�B�R�CMQP*��b !GCLF�#�1DY�8} �q�35T�%DG���0��5I��SSt0��BC P��1�A��`Q_�1�8�11��E�C��13 K5 F�GR)A��gC��k�`�W�ON��"EBUGwctBx��C ��_E D ����` �TER�M�EE�EA��OR�IS�@F�E���S#M_�`���@G�E���TA�IH�E� I��UP��I� -�Q��D|`�C|P�E$SEG#Z�0E�L�eUSE�PNFIzLRT�kA,��D�TF$UF�`O�C$\��a�P/��ďWi@T��t �cNSTTPAT��h��ROPTHJKa-�E
� 65MR<p&�WUw�&�Q��LQR<`�Y�qSHF�T��MQ�Q�X_SH�OR�*��F �@$��GM`H�u OVRHq��q6`I`4U�= �aAYLO���"J�Iu2b��Q��oƸ�ERV���a� 6j� �WnP�R~�E �e��E �Rb1Pp�ASYM|�p�MQWJ`W�� AE���Qy�b0�U7t@nPI��Uw�/�ePo�X�`o�fgORnPM��G@SMTfJ�g�GR��aC�qPA�|P���=��K �� FTOC�FQ�P9`N $O�P@/��#��N ��!O�ڐRE
�R�dS�QO����Re��R�UN�%�a#eo$PWR0IM@���bR_ �L�=�mR �LVBH�_A�DDR$�H_LE�NG�Rǁ���T�R�� SO�M H�S ���~��������	�SE!u���HS�:�MN�1N���p��F¹�OL���8�3�3�=��ACROc�z�P$��[�p�a;�  �OUP����r_�I���q�q1 �ѭʓ��ԙX!՘Y1 ՘t!՘	�ԙлE"IO���DϗA�ߕ<9�gO $���p�)_OFFb�;�P�RM_Ò�1HT�TP_[�HjP (��OBJ�2��#[$$�LE�S��>�Q � ����AB_�!T���S��p;x LV��KR�32@�HITCOU�BGE�LOہ 磴!��@��"�G#�3SS��HWD�SQ�jR�lpINC�PU4BVISIO �����Ğ�
������~	� �IOLN�S� 0C$�SL�r@PUTM_�$@��PV0x�ɱ)F_AS�2T $L  �� D=a0U�@9`dQٵ��䳊`HY#�]�6Ù���UO�3U `"�{�$�5"M�5 Tƥ�R�P;@��ǿ��T��µ��AUJeV�]���NEfgJOG�{W��DIS���K���� �3W XХQV8v��P;�CTR�S:��FLAGBB��LG�tX �� ���aC?LG_SIZ���`��d �����FD��I�اؓ�׏ث@�� �����	�d 	��	���	�@	�% SCHA_��R���aBg�N�*��Y��!E�2��p�J U}�}��pL܆�|�DAU��EA`�����t���GH�r��%�BOOZ�h A<�f0ITp2���@8�REC�GSCRB�=�D:�<����MARG�<1�8��0��a�%�S�ȣ$�W?�%���0�J{GM��MNCHz�%�FNKEY��Kn��PRG��UF���g`��FWD��HL.	STP��V��mPX������RS;	Hp��-�Cid6r0�.0s��	U|���r�Xb���P�E���G��`PO��
.�M�FO{CU�RGEX,ǗTUI��I��p� K|�V��V����A`@B���p�A`�Nu���SANA%�FR��V7AILy�CLP1u?DCS_HIyD�D
��O�X1�S� ���S�V�IGN ��~�ӽ�\�T���^%�BUFF�1[5�5o`T�$��� H����B�f�A��\5�o`ܰ��c��pWOS1�%2�%3�!�P$��0] � �ܩ�qEU�����IKDX�tP�bD�O� X��Q6ST|�R���YV�@1 \$EO6CO;�{�^6q6q�$.��1^ L�� K�[@`�9`(��S����:������%�_ _ �pp�Ð���t C�@Cp�` �� �CLDP|�uTRQLI��Ft
�4I"DFLGV�"@1VC�1D)�VGr�LDVE@DVEORG
�qiB_瀶g�H
��d�D�ta� �M�@Dr1DVESB�pT4@I��@TVRCLMC%T�O�O�7Y���MI��tb� dy��!RQI��M�DSTB�0 ��VO�XAXr ��X�\EXCESH6���vRM_��qc6���Rt�1vR<��pd��V_A�Z��(k�_�X@K�te \�����/�$MBs�L�I���cREQUI�R�b��l���hDESBU��sQL�0M,Ձf�r=��`����%RFsQND���p�pgw�n�?�sDC��I�N����p�,x' NpV���K�NV�cwPST� h��7LOC�&RI���%EX�vÀ�!�QsQ�ODAQ,�i Xf��ON���MF\� ���v9�2%��5�uk��0� �FX�PIG}G�� j �M�@�2!���3��4R �%?3;�|�K�|�Z�<G`E�DATA{'��AE�U��b"���NZ"�k t $MD
��I��)Ɔ ф��фH�p�`Ѕ�X�҃ANSWe�ф�!'jхD[�)��MO���P��l �PCU��V�X@�uRR2��m D���a���R?d$CALI�P"��G�w�2��RIN���z�<P INTEڰ�"nI���°r��ڰ_N��oÕޒi��oT۔bp�DIVFmVDH�Pݐ��q� �$V��+s1$��$Z�"��� �"�f�_�e�rH ?�$BELT>��1_ACCEL!������IRC��P���t�T31h�$PS�P'BL��M�ʤ<Cඐ�������PAT!H������3ТZ��Q_�!U�2�8�R� �C堌�_MGP��$DDU���/�$FWh�����q������f�DE��PPAB�NاROTSPE!EH��!��4@J��!���P����$US�E_���P��O�S�Y��g�Q B�YNryPAO��OFF�n�MOUR�NG��O�OL�L�INC .��q��u��Rn�PP�RENCS�����RȡX���TŠIN'2IТ0���`R�VES�{�>��23_UPI���/LOWL!� �4@���D� �R{`����0��5bCΐ��MOS4 LdMO���PWPERCH   �OV��b��!m�@1 �^T@1�s��hP�`Ä� V5�'`ѡ��L`���Ig����UP��8����TRKv�#2AYLOAA��$a�1�Т@�5�p40��RcTI(a|�40MO�� ��R$b�@N��T��w��L���"f�DUM�2,�S_BCKLSH_CТ��B�A� u�'�Y������6�x�aQCLALz ���A8r�`�CHK4@+5SH�RTYS���}%�A��_:36�_U�M(`n�C{�c�SC�L��ʰLMT_J'1_LS��P������E�����������SPC��;���	&��PCsѦ�H�0�`dY�q�C3P�2XTc�.g�CN_��N��i"��SH ���V	�*3@�Ň�=Т�AC� y�SH:3��g��ƝA ���s�4�ѡ��c�3PAx�l�_Pw�[�_5@��8�V�4AH�Z�K�JGG"M��OG|[��TORQU��ON.�Q靰wbLҠ�L���_W��1�_A���G��M��I�IJ�IM�F�p�JPQX2(�A_�VC��0�T�RS"1Y.�Pm/�R`%�JRKY,�"�&PD�BL_SMh�RM�)p_DLG�RGR�V��$G��$M��!H�_ �#�:COS;`�8LN� ;;\% B4G�=9M�=9!y:g<�-!�%Z60L־!MY�D1�8$2TH*=�9T�HET0�NK2a3M�BA�E0CBFCBA�C�Q�R,B$0:AG�:AFSBG�XBNEGTSaʱC� �qW4&�Dg3�Gv3$DUH�Ih�Aw� x��R�F���QQ���v'$NEd�IF0Y�H`R�E��$%��1A�5�#U,W
581LPH(eR��RS\%tSg5 tSv5R�6�S�Z�6%�EVEXV:X7�]\VlZUVy[V�[V�[V�[V�[V�YHEX^VdbP\]�{hy[H�[H�[UH�[H�[H�YO6\�OEXO�i[^OlZO�y[O�[O�[O�[O
�[O�6FR'A�yg5��t8WSPBALA�NCE_�1�sLE6o@H_�5SP��X6��rg6�rv6PFUL�C�x��w�v5Ț1=n}�UTO_C�n�T1T2G���2N *�z���g���k���@(ע����T��O���>�INSEGz�%��REV��%���DI�F��1o҇�1p�@OBȁ��#���MI��5��$LCHgWAR����AB*~y�$MECH0A��0>�D�Y�AX>�P���]�W(�<�q 
p^������ROBVУCR�Ҡ�R��M�SK_�pj�s P+ R�_��R��H�Ҕ��1���ԲҐ�����Ґ&�IN����MTCOM_C|D n�t  P��ڀ��$NORE���9���(�u �8�GR�I�SD��@ABJ�$XY�Z_DA9Q���D�EBU��M��U�vu �p$�COD��G ��o�J�j��$BUFIND�X԰����MOR^œw $1�U�� -��v�F����Д���Gܢx � $SIMULX���x��$���OBJE�p>$�ADJUSB�5�OAY_Io��Dc�����G�_FIJ�=�T����������������Հ�P��DN�FRI��׵T��RO���E������OPWO� ɐy�0��SYSBU<�PΠ$SOP����#�'�U&�ՀPRUYN�M�PA�DLƸH�!���_OU�!�A���r�$��IMKAG��ϐ�@P��3IM����IN� u�~��RGOVRḎ>°Ѐ�P����԰�@�L_:����m� R)B� �@M��SEDՠJ� ��Np�M.���^����SL��pɐz x $�OVSL��SDI��DEXqk�i�=!H{��Ѕ�V���N�р�{��Њӟךط�Mx�!РF�_SET�ɐ{ @���g���SRI&���
��_4A���	����ׁ@��  �| HϑI�J�A�TUS��$TR�C�@ǰˢD�BTMTM�7�Ij���4��#�,�ɐ} DϐE~�k�A�`EۂBᏱ8
��B�EXEH�Z� ќ��{���~��АfG�UP���$����XNNm�=!p�L!�p� �PG&��!UB6�g��6�~
�JMPWAI� �P��N�LO��j�F���#�$RCVFAIL_C�j�Q�R��Q�Z�M� 𣕠����0R_PL
�D�BTBm�j�BW�D��A�UM���I�Ge���m�� TNL�� ����R���.�E�p���DEF�SPy� � L�ϐd�7 _: H�HUCNI��r�F ��R��,^�� _L��P@�0 ��ȑ����F�����Ѐ��p��N�pKE)T�}�� P��ȑ�� hW�ARSI�ZE��l���S�@�OR
�FORM3AT3���COJ�����EMV�lU1X��ҎLI��ȑ��  $#�PO_SWI�i�G���AX����AL_ S��E A��B��,@C��Dj�$E6���uC_��	� � � ����qJ3�@����TWIA4�5�6��MOM������4�#�Be�AD�&��&�PU;@NR �J%�J%��HŔ��� A$PI �F�ޑ��$�%�#�% �#�%=D�&�+QD�Dpф�F���U���g�S/PEED�`Gd*4 f�7167f���16�g3@8��O9��f�SA�M�p맣417�3f�MOV���D�1ƀ�E�4H�E�17 1��42�@������5n��Hm��3IN2Ln�39HUK�0Df�;J{HRD{K�KG�AMM�v�A�$GGET��ȠL�D�z �
b�LIBR��I��$HI��_���P��bVE�XA^:P+VLW]XVO\ :Y|V+V�V������ $PDCK�U�L�_�0�� �.B�m!E�W��T�&�Yr �$I�RS�D��&�����(�LE�ޑ�OhĤ)`�s&�ɐ��P��UR_SCR���a^��S_SA�VE_D�īe��NO�C����`�D ��&�i��)�iapz {p���&Ex@�q� �0�B���5G�2�+8 !�;6��g8�w�ucs�1���FM{%� ����!G����c�w���`ζ�qW�`��$���0�N ��R�qML��H�CLG�GM�a�ǒ� � $P9Yr�$Ww�+�NGt��w��u�� u��u��������@([L�nX� O�m�Z��GQ�Ŕ� pW�#�c�&�o�o�#5��_)�� |Wи�`������@��`�ޗɖ�EQ�P�Eg���b�Ϡ����P��PM��Q}U�0 � 8� �QCOUas�QT�H��HOL��QH�YSES�1[�U�EG��b� OM� � �P4�U�UN\I�J� �O��)�� P�������a��ROG�j��2��O𤥥c�󠉠�INFO(�� Ж�ث�
�ȏOI��� (`SLEQ"6D�5D�ܦ����IDS𿠒��VPO�P��0#3QEMPNU�����AUT�a��COPY�1�಼��`EM��N������CT��� �RGADJ�(���X#�_$P� '��'�W%�P%�`]`'�:3�;�EX��KYC���@OՐr(��BЗ�_NA�1!S���i����M?� � ��p��POR��Ì&��S�RV��)����DIT_p��� ��
�P�
�w�
�5�6�%7�8��1S�b��=���MC_Fe���pL�a�a�;�R q���/��җ#�0���k��� ,`FL�����`YN{���Mzp�C��PWR��������DELA4 �6Y�ADR��� �QSKIP{%�� �����OŀNeT�1�0*�P_�� ��I�`߂̐`��#`� 3`��n�kn�;�m�@H�m�U�m�b�m�98a��J2R.0��� m4� EX�@TQ� ���q����������jRDCx�� )���X��RF�E�@AY�_�X�DRGE7AR_�@IO�t=b�FL��Q��EP9C��UM_���?J2TH2N�# �O 1�UA�G�@�T�P �"���M���-�I���4?�EuF�11(�� l!��ENAB� ��TPE2`{� 8Wܠ �M�q�CL��R��w U2'� -?Qcu���3'������� S4'��'9K]o�5'�������
6'�!/3/E/W/(i/{/7'��/�/@�/�/�/�/�p8'�?-???Q?c?u?�SMSK(������ E�aM�OTE���
�`�`/B`��q-CIO�U�QEI�0�p&�R� W\`��� /���-�����ҿ���ՈB$�DSB_SIGN�'a�q����C��pE^S2323E����$�DEVICEU�SKC�r�rPARI�T!�AOPBIT��q��OWCON�TR���q�0�rC�UPM�sUXTA�SK�SNq��P�DT�ATU�p)BS�3`���u�e�_�pC���$FREEF�ROMS������GsETA`��UPD��9AEbxaRSPTP��߫� !�8$USA�����9h�{��ERIO���`ՐRIY�U�B_�`�P�Q�QfWRK�?�<D�h�3fh��6FRIE�ND�qg�$UFx�U�p`TOOLwf�MYd�$LEN�GTH_VTߤFcIR��cM�SE�@��iUFINtrа�ARGIaF�AITIi�gXF�i�fG2�WG1�� �S�r$wPR��sau�Oa_�@�P��xQRE��0�SU�ءTC�N�=qyv �G��]R���u��Q�A��hzh ZUz�ZU�t���{P�T��X �P��L
��TcH��hh�U��T�SG��WX�)��r>�D���.��C�z�N�b��$�v �2�!�-a' 3i1T?h.`21k2��31k3?j���@i����60{��s{��r$V��b�V�eV���vYr���O�[V{�@��hv3R0u�^pib��PS���@�0��c�5$A8й�PR)��u,�qS���@���U��¯ 0p�v���P�N����!��P>p 갢
�USzA� E�\�R��GA_�Š���Ny@AXQ��A�g`L�ag�p�THI�C'a��-����QT�FE���m�IF_CH'cp�I_����6D�G1՘٤*��h��`��_JF�P�RW�I��RVATF�� �\�'�f`���)�DO�e)�CO9UW�C�AXI�D��OFFSEZ�TRIG�sz�,�)�#g����z�H����g�IGGMA�P�a\����ȸORG_UNE9V#@Ͳ �SD��?�d �$��=��GROU[A��TOa�Q�DSP�#�JOGV�S8�_	PV�3RO���U�mpnEVKEP��IR?�d_�=pM ���AP����E�������SY�Sv��B��PG��B�RKYr����b�\�`�������k�ADVQ<�y�BSOC�C@�N�DUMMY1�4��`SV�DE�_OP1SSFSP_D_OVR�� 1C~�N�Q�OR\׶0�N�P]�F��]�<�OV?�SF��a����F���Ac�As�؁a�B�LCHDL�REGCOVM��P<�W�`1M<��?�RO1S�rK�_a�_� @����`VERt�$O�FS�`CV�@_bWDv� �r���R��9��TR%QA�E_�FDO��MB_CiM[A��B/�BLl�_¦�l��V�qDb�PȢ���G���AM��Ú�yP��'��_M��>R��HC4�8$C�A2���Ȱ��8$HcBK�Q��N�IO1eq]�iAA�PPAQ��}�b���u��iB4�DVC_DB�c�� �B����A��1��'����3��-�ATIO"�@��FPM�UDc1�HFCABH�0bFs�p �p��Ea<�_BP��?SUBCPUk�I�S%��@����P�s��,���B��$HW�_C!��i��x�A�'q\�l$UNIT��l�AT}�����I�CYCL��NE�CA#��FLTR_2_FIҤ�H)��FEaLPU˲���_�SCTosF_�F0��
v�
FS�A���CHAJa^���3R�RSD1�B �ؑ�l�i@_T��PR�O ~�)PEM�0_����8�3� ��<�*%DI�P��R�AILAC��rM���LOГc+�i�`��-��-'�PR��%S{q*��!C���@=	&�FUNC�³�RIN�pZ�+`? �$f(QRA� mr 9�p�#��G��#WAR�F:�BLuq�'4A;88DA���!I835LD�PA�A�q3dh��!��q3TI��p�5�β�pRIA�Q�BAF� P�A���1@��5��T���EMJ�9I1Q��DF_�`��l�Q��LMt�FA�`OHRDYd�P�`�RSoq+`Q0EMU�LSE�`���E�G ���I������$]a$�Q$�Q�,��� x��EG���A�ƠAAR�2)�09pmb�E50��AXE&ǗROB#�W�ac�_�M�SY���Ae�VMSWWRذ�M12�� STR"Ņ�d�h�E� 	CUq#��lqBhP3�oV��)��kOT�P� 	$�ARYg��R_!�`�	T�FI��j�$�LINK�1w��Q��_eS3�CU��RXYZQ��[��	c�o��Q�R�X�PB!��"Kd�
 � LcFIeg3�D�9Ԫ$<�_JN�"�e��SA�'OP_~T�[53�Nq#TB�aNB�bC9���DUQ�BV6r%TURNb���u�Q�!h�?�gFL)���B�@�+pekZ73�I� +1�nPKH�M��BV�8r%����c�ORQ&�!�#mX�C���� �갦��u��.�<��t'OVE�q��Mj�@tC�zC��B�W� Fq�� ���� j�0 ���qw�P����	��q����zC��5��!ERM��!	v"E8P���#؄A����id�%"�WP1MP1AX�bP1 ��&!�Q2�2!>�\A>� ��=��`=�p=�ep=� �p=��@=�JQ=�@:� @J�@Z�@j�@z� @��@��@��@���ב˙DEBU�$�!�1(${�P��R�g� � ABP'N�[��s9Vְ� 
���� ��Ϥ��Ϥaڧ$aڧ �aڧqڧeqڧ�qڧ��A�4�`�2�RLcLABbb�u� ���1so 	�ER�>9P � $8`� mA�!��POB��FЉ�P����_MR}A��� d O09T<�\�ERR:�2��0TY�aIA�V8b`,���TOQ+�i�L�@,�7R��p³�о�A � p�T8�P��< _V1ْ.�(V�2#c�2\�2k�ȱ���op�ˠȱu�$QW��6�V�A���$�"�0,���6��Q�	�@HELL_�CFG�A� }5e B_BAS���SR��p�� ��CS��1�1��%��22�32�42�5*2�62�72�82���RO �8��P,`NL�zA�cAB��H �ACK��>�i���`�`�G@���_PUr�CYO�@��OU��P0��W!��3�7LTPX�_KAR���RE��&@P W1�QUE� �p9C�CSTOPI_AL�����Pq�Д�ఎ�PSEM���Ml���TY��SO��W�DI����}�L��1_TM�MAN�RQ��PEZV��$KEYSWIT�CHq8��CHE�9BEAT!�EF�@LE�$f�U4��F��5�K��O_H�OM�0O�#REF�pPR�!)�AUP���C��Op�0ECO�ư_1`_IOCM�d��������g��@� D�Q� U�۲{�Mw2Q��p�cF�ORC�3 �5���OM�@ �� @���3�U[SP��@1��$�@3�4��1[NPX_AS��¼ 0�ADD|' h�$SIZ�$VAR2�D@TKIP���� Ah�аJ�� �� �B�S��AC��%FRIFa��Se�w	��NF�@Џ@�� x�SI�TE�Fsj"esSGL}T�R7p&A���#P~OSTMTJ�P�@�;VBW�pSHO9W�R��SV
@�D߿� �ԱA005pЁ "� '� 'P� '� '5)6)U7)8)9)A) �@'v 'V�	&r`'F(JP�()�P�(,) #`�(F)p�(`)�p�(�z)1�)1�)1�)1��)1�)1�)2)2�)2)2,)29)2�F)2S)2`)2m)2�z)2�)2�)2�)2��)2�)2�)3)3�)3)3,)39)3�F)3S)3`)3m)3�z)3�)3�)3�)3��)3�)3�)4uI4�)4)4,)49)4�F)4S)4`)4m)4�z)4�)4�)4�)4��)4�)4�)5uI5�)5)5,)59)5�F)5S)5`)5m)5�z)5�)5�)5�)5��)5�)5�)6uI6�)6)6,)69)6�F)6S)6`)6m)6�z)6�)6�)6�)6��)6�)6�)7uI7�)7)7,)79)7�F)7S)7`)7m)7�z)7�)7�)7�)7��)7�)7�$5�V�Pd�UPD�� � ���)и�Y�SLO��� � ����Q��T�A�����ALU������CUT��F���ID_L��H�I�IV$FILcE_�?�+�$��v��SA��� hҰ~k�E_BLCKh��x����D_CPU ��� ��� �B�T����q�	�R �G�
�PWl�� �L�A1S������RUNu������8��u�?���?�� �T�?�ACC���X -$f�LEN@��s���f�����I��J�LOW_AXI�h�F1f�,�2��M ��	�G�_��I��Y�8�թTORn�f���D��ܣ\LACE���Y�f�ٳY��_M�A� ��3�	�3�TCV:�[�	�T�\�{��q�|������	���J$����MĴ�J9��R���	�r�2��`��������ΠJK�CVK��#���#�3óJ08�'�JJ/�JJ7�AAL'�]�/Ô]�W�4X�5��{�NA1����M�I�ڤLӠ�_���b����{ `u�GROU�����Bd NFLI�C��REQUI;RE��EBU��b�Ŷ��2�c�	�xa�� �� \/APPR�C �ܠ�
a�EN\�CLO��l�S_M`�������
a��� �F MC6�{�����_MGV��C�l��ظ��5���BRK��N�OL�����R�_CLI�������J��P_��/��7��{�����6L�O��8�[b�?���# ҍ�z��燡��PATH�������ᒨ��� $��ͰCN��CA �]���INe�UC٠��%�-C��UM.�Y��4��Ez�P���P�7�~PAYLOA��J2L��R_ANE���L����������R_F2LSHRC��LO��$����2���2�ACRL_@�"� �����H��b�$H��CFL�EX_�`�Je�� :r���	�t������	�������F1���ïկ�����E'�9�K�]� o����������$�� г�#(ؿ�����TR'�X ˲� `H��%�&�8�J� \�`�i�W�{ńϖϨ���_��� �� ������ʁ��A�T�ðELt ��5�J����J�E��CTR�T�N"F�6	�HAN/D_VB�_��n��� $f F2�����SWF������ $$M����R�ӅH�ѕL��E:�FA�������I���A��݀��A��A�	��@�۪���D��D�	�P��G	�qYST���yQ��yQN�DY  �Z��ּD�E��)��� �������H$� � �PT�]�f�o�x������J>�� �{@`��n�vf��o�A'SYM�������Ͱ����_SH ��#�=�'��dLHG�Y�k�}���J��G��gs�]y��_VI/C��x�ӵpV_UNI���t�#��J��re �r���t���t�ð@	G�(:j��#P�X}1A�H��N���EB��EN/@��DiI	�W#O���`������� � �BI�aAK����吂���U��0`��n�� �[ ]AME\?0h�g���T��PTp i0��5�����K�,p�:�U�I�TKp�� �$DUMMY1��!$PS_RMF�   ����͑LA��YPV#��=�$GLB_T~@ ��ŕ5���`�CAӁ�� XI�	נ�ST�ȱ�SBR��M�21_Vɲ8$S/V_ER��O���#�CLߐ�AuO�炔��0O� �o D ĐOB���3LO�f�S�y�Ð�S�p�1SYSS�A�DR�1��5�TCH>�@ � ,f L����W_NA
������1��SR>��l }J�J ���F��B���G���I ���ID���D���D��� V�p�KYV���bu��� ݻ������);Mt>��XSCREi�W�5�E@�ST��F��}��a�Ǥ����0_�0AV�� T I�&����1%�������1�����O�PI�S�1��� w�UEЄ� ��䪠��SG��1RSM�_����UNEXCcEP��ј�S_ߑ ��7��&�9�T����COU\ғ� [1֤�UE��؂|6�y�PROGM@{FL�1$CU&��PO�>��UI_��H�� � 8\E��_HE_�������RY ?��0���������OU}S � @��~D�$BUTT/��R����COLUMx0��s�SERV�3���PANE�0V��:�TpGEUA|��F��ʡ)$HELyP��bETER5�)��E���Oq��30�� ;0��M`��U`��]`��SIN��-�TpNp���0�131� ��i�LN��ܓ �0���_����s$H_�0TEX�3�j�^�~$RELVB"D��~Ӑ�b���Ms�?,��p��4������#��USRVwIEWV�� <����U"�]@NFI<�0��FOCUA���7PRI�`m��h�� TRIP��m��UN��Є� x�`/��WARN�����SRTOL���&�Rs�O�cOR�NsRAUW�vT��	���VI�υ�� $��PA�TH���CACH�V#LOG��LI�M�r�S��BR'HwOSTǢ!�z��R|�OBOTƣV#IM� ��S����0r�������V�CPU_AVAIYL���EX�!�aN��} ~�Ma�Ua��]a ������$BACKLAS�� �!�$"W��  �CT%s�@$T�OOLǤ$�_J;MP�� ����$SS�v4��V�SHIF`у�APB���ǤЇ�Rk(^�OSUR�3WRADI�$��_ ���%�м1�ぺ��$�LU�q$OUT?PUT_BM��IM���b� }p���#wTIL�'SCO�"�#C���$N�&N�' N6N7N#8����u%=,�2����V��υ�<��D�JUrU��P�WA�IT���<��:%�0NE~��YBO�W� �� �$������SB"IT;PEo�NEC/,B@@D(D�PJǐp�Rv @hE(�#=@�0�B�E/�M�KT���"y�� �An�!�OP�
MA]S��_DOآ�qT��D]����C��>RDELAY��SJO�"X֡�c'T�3���`� ��,l�y�Y_Ry�wR�#Ƣ�A�? ɀZwABC�� ���R��
  ��$$C�X�����Q���P�P�PV�IRT�_�PAB�S�!��1 �U�� < �Q(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�K�|`�AXLMTZvK��c  �]��INf�x�\�PREȏNk�����LA�RMRECOV ��Y�����@F ��U�QdK��"�4�F�T����w���������,c 
#o�W�NGu� k	 A �  �,�`PPL�ICu�?�U����Hand�lingTool� m� 
V7.?70P/36+��;
��_SWr��F0���� 43�ˊ�yϋ�7DA�7�철
f��{rm�None�����Oհ�P�T_���<�_+��V��R�v�7�UT�O�RX l���n�HGAPON�Pe� an�U' D 1�� �и�����T�n�ދ Q 1�  T��������	7�0H嵡]��R�P�Qg�a�,�H����B�HTTHKYV��R�+�=�O�� ����3����!�?�E� W�i�{����������� /��;ASe w�����+� 7=Oas� ����'/�// 3/9/K/]/o/�/�/�/ �/�/#?�/�/?/?5? G?Y?k?}?�?�?�?�? O�?�?O+O1OCOUO gOyO�O�O�O�O_�O �O	_'_-_?_Q_c_u_ �_�_�_�_o�_�_o #o)o;oMo_oqo�o�o �o�o�o�o% 7I[m��� �����!�[����TO�C�U�DO_CLEAN��5Ի�_NM  	�Կ���+�=�O���_D?SPDRYR��HIa��@����ϟ ����)�;�M�_�pq�������MAX@� ��[����׳�X������҂�7�PLUGGp�У���S�PRCt�B���������O�}�5�SEGF{�KY�k�v�������Ͽ���=�p�LAP����o�Y�k�}Ϗ� �ϳ�����������|1�v�TOTALզ|��v�USENU����� ���ߎ���R�G_STRING� 1s�
�kMl�S3�
�ѿ_ITEM1��  n3������"�4� F�X�j�|��������������0�B��I/O SIG�NAL��Tr�yout Mod�e��Inp��S�imulated���Out���OVERR�� =� 100��In� cycl�����Prog Abo�r����~�Sta�tus��	Hea�rtbeat��MH FaulAler%	U�C Ugy������ ���۞��� �6HZl~�� �����/ /2/�D/V/h/z/�WOR y��۲!&�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO0NPO��V@�+ ?OyO�O�O�O�O�O�O �O	__-_?_Q_c_u_��_�_�_�_�_QBDEVYN�PmO�_!o3oEo Woio{o�o�o�o�o�o �o�o/ASe>wPALT�q �/x����� � 2�D�V�h�z��������ԏ���
��GRI����B���j�|� ������ğ֟���� �0�B�T�f�x�������0�j�R�Z��� � �2�D�V�h�z��� ����¿Կ���
���.�@�R�ԯPREG �~����dϲ������� ����0�B�T�f�x� �ߜ߮���������X���$ARG_� D ?	���9���  �	$X�	[�M�]M��X�n�,�S�BN_CONFIOG 9�������CII_SA_VE  X������,�TCELLSETUP 9��%  OME_I�OX�X�%MOV�_H����REP��S�&�UTOBA�CK�����FRA:\x�c Z�x���'`��qxǣ�l�INI�p�x���l�MESSAG������A�>��ODE_D���ă�#O�P2l�PA�USVA!�9� ((O<��� ����� (^L�p��e~j@TSK  ux����o�UPDT) ���d ?WSMg_CF��8����%�+!GRP 2
V5+ L�B��A��#�XSCRD/!1�5+ ����� ��/�/�/??(?�� ���/p?�?�?�?�?�? 5?�?Y?O$O6OHOZO�lO�?O(�r�GRO�UN S�CUP_kNA�8�	r�n�F_ED��15+�
 �%-BCKEDT-�O0�%_LI_�� ���-r�_x�o�o�x���U2r_/��_�_�R��o�iU�_&o�_�_ED3o�_�o�_n_o8�o9oKoED4�oro�'�onn�o�oED5^�:n�8���ED6���o��nK���%�7�ED7��^����n�8Z�ɏۏED8J�*_��N_m����m���ED9�[�ʟ`m7����#�CR_ ����7�ٯD���ū��@�@NO_DEL��O�BGE_UNU�SE�O�DLAL_?OUT ��R��AWD_ABOR��𦾦AݰITR_�RTN����NO�NSi ����C�AM_PARAM� 19�#
 8�
SONY X�C-56 234�567890H ���@���?}��( АZʨ��yŀ��\�H�R5o�������R5y7����Aff�� \�L�^�Z��ߔ�o߸� �ߥ��� ���$�6���Z�l�a�CE_RIWA_I(%;��F�!{�x� ��_LIS$�c%����@<��F@�G�P 1Ż����OK�]�o�.�Cg*  ����C1��9��@��G���CVP C]��d��l��Es��R������[��Um��v�������_�� C���& ���G��;�HEנO�NFI���@G_�PRI 1Ż ��T�������� �CHKPA�US� 1I� ,�BTfx� ������//�,/>/P/b/t/�/Oƭ����8�!_MkOR��� ��@�#B�*���% 	 �)?�/(?? L?^;�"����-=�ֱ?99��3�@K(�4��<P������a�-8��?OO�J
�?KO�'ưS����:O��i`��P�DB� �-+�)
�mc:cpmid�bg�Od��C:� � =P>���Ep��O-_�C  �"������!S�@�O�q_<Z�  pPqS[_�_=Y�*,��,��S[g�_oV�\�װ�S[f�_�KoAMo�JDEF 3ch�)�B:`buf.txtqo��Mro�0����'�	z�A��1=L���j+MC�#�-,���(>ss�$�-�r���Cz  BHF3C�s7 C���C��M�F��iDP�E�~�WJ�I0D�tE�q�aEpIJ$��3HHƷ���{F��G���GG���N�[5K~w)L���XWI���fu7���4�)�.װ��,�,��@�u�K�)x6�q�* �* e�3D�n��pEWLI0�EX�EQ��EJP F�E��F� G���~^F E�� �FB� H,- �Ge��H3Y���z�  >�33� ���|F  in6�|A@��5Y���<2��A�1WDq<#�
 �O+�)�Zj~�bRSMOFS����n6��iT1� D�E  �?DR 
��,�;�&�  x@�:��nTEST�b)o�8�R��!�/3��nvC+�A�WJq� �[��rq�C�pB�1 w�Cy�@T�6���T�FPROG� %ź��ů��I����𦶠喤KEY?_TBL  �6Q��!� �	
��� !"#$%�&'()*+,-�./01g�:;<=>?@ABC�`�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~��������������������������������������������������������������������������������������������������������������������������������������������L�CK�X	���ST�AT*��_AUT/O_DO���G_��INDT_ENB�K��"R��i�[�T2<��\STOP���"�TRL��LETE�����_SCRE�EN "��kcsc��U��MMENU 1""�?  <���� |�WE[߅ߺ�V��߽� ������,���b�9� K�q��������� �����%�^�5�G��� k�}����������� ��H1~Ug� ������2	 AzQc��� ����.///d/ ;/M/�/q/�/�/�/�/ �/?�/?N?%?7?]? �?m??�?�?�?O�? �?OJO!O3O�OWi;�_MANUAL��ޞ�DBCO��RI�G�4�DBNUM��`�<q*�
�AP�XWORK 1#"�ޟ+_=_L�^_p_܂[�ATB_�� �$"��ipT�A_A�WAY�C
�GC�P *�=���V_A!L�@M��R�BY���4*��H_�` 1����_ , 
^7��6�Boo�f�PM��I�j��\@��cONT�IM��*���fi
�$cMOT�NEND�#dRECORD 1+"�qer9�a�O�Oq =6��R{���Hx ��O�s(�:�L� ��������ʏ܏ � ���$���H���l� ~������Ɵ5��Y� � �2�D���h�ן�� ����¯ԯ�U�
�y� ���R�d�v������� ���?�����*ϙ� N�9�Gτϧ`�^�ϼ� ��=�������(ߗϩ� ^�p��ϔ�����9� K� ���!�H��l� ���ߢ��K�a���Y� �}��D�V�h���R�TOLERENC��TB�b�PL����@CS_CFG �,0k�gdM�C:\��L%04�d.CSVi��Pcl���cA CH z�Poo�n"W^m��c��RC_OUT -�[=`�o��?SGN .�Ur��Q25-MA�Y-20 11:�00 ��af P�X��n� ��#�pa��m��PJP��{VERSI�ON �
V2.0.11�k�EFLOGIC {1/�[ 	tH��P��P��PR?OG_ENB�_r��ULS�g �V��_WRSTJN�`�F��MO_O�PT_SL ?	��Uac
 	Rg575�cO 74T)56U(7U'50y(t�"2U$tH�/z2$TO  >-�/{[V_�`EX�Gdu�3PATH A�
A\�/]?o?��kICT	aF�P�00g�Tdc�eg��1STBF_TTS�h�I�3U��Cda�6�@MAU� ��bMSW��1D0i��l� ��2�Z!�mO|3bO�O�O�O�O�O�O_tSBL__FAUL� 3�_|�cQGPMSK�^�bTDIA��4�=�d`��a1�234567890�Wc|6P�/�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o\SZpPf_ *��O R*�?%�PBhz� ������
���.�@�R�d�v�H|��U3MP4!Y )^���TRNBKS��ĀPM�E�5ЏY_TEM=P��È�3��D3�����UNI.��Y�N_BRK 5�����EMGDI_�STA%�W�NC�2_SCR 6G��_����͟ߟ�f ����0�B���~�e�17��;������¯�,R|�d�8G�� a�������N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶�0������@$<� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ��������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/� �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gO�/�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo�Oqo�o�o �o�o�o�o�o% 7I[m��� �����!�[oE� W�i�{�������ÏՏ �����/�A�S�e��w���������קETMODE 197��v� '��� �W�RROR_PROG %��%���X�'�TAB_LE  �A�𚯬���њRRSE�V_NUM ��?  ����)�_AUTO_ENB  #��j�w_NO� :��
��  *�*F��F��F��F����+E�_�q����HI�S�h���_AL�M 1;� �2��F�F�+�� �@�$�6�H�Zψ�_�.%�  �D�����ېTCP_VE/R !�!F�j��$EXTLOG_7REQ�������SIZ����TOL�  h�Dz����A ��_BWD��5��a�	�_DInO� <7���	�h��k�STEP�w߉�ې��OP_D�O��4�(�FAC�TORY_TUN���d��EATUROE =7�a���Handl�ingTool �7� DER �English �Dictiona�ry=�7 (RAA VisS� Master0��>�
TEa�nalog I/O7��>�p1
a�ut�o Softwa�re Updat�e�� "`��ma�tic Back�up;�d
!���ground� Edits�  �25LCa�mera��F�� w"Lo��ell���>�L, P��om�mj�sh�8�h6�00%�co����u�ct%���pane�6� DIFD�'�t�yle sele�ct�- `�Co�n��j�onitoir<�B�H��tr5�?Reliab�� ��(R-Diagnos���:�y��Dual Che�ck Safet�y UIF��En�hanced Rob Serv��q (V�U?ser Fr����T_iE�xt. oDIO ��fi��u Z�\=end �Err��L��  �pr�[r��C  �P���ENFCTN Menu��v����.fd� T�P Inp�fac��  
v�G��p�l�k Exc	 g�5t��High-wSpe Ski��_  Par\�H��~G mmunic��wons��\ap�ur� p���t\h�8��con�n��2� !D�Iwncr� strZ��i�<�M-6< KA�REL Cmd. L� ua���8~sRun-Ti4 Env=�(mqz �m�+��s��S/W�=�"y�Lic�ense��' a����ogBook7(Syo�m):���"MACRO�s,�/Offs%e��f���HG R����M1?�Mech�Stop Proyt��d 5
$�{MieShif���9�B6SD�Mix� ���7�y�Mod�e Switch���Mo����.& R�M�&��g' 6�5�ulti-Tp� ����Z�Pos���Regio�  �! 7Pr�t F�unb>�6iB/1��Num ��d�x�P`�312  Ad�ju:�/2HS�M7Z* oY�i8tastu1<�AD �RDMotN�socoveW� #���3�uest_ 867.�9oG �� �SNPX b����Z#Libr<V�;�rt IE,�� S$@�.�0�� ��s in VC�CM9��0�� `��!9�3��/I�� 710< TMILIB�MJ0,@� ��Acc����C/2�@�TPTX"+QTeln �Lq3�%�|(PCUne�xcept motn�� �0�0,	7�?\m72f�+�4�f�K  h6�4aVSP CSX�C9�@(P�U["3� 7RIN�We'g50,D��Rvr��	menS@� �Qi�P^ a0��3fG�rid�1play F O`�fp@���vVM-�@A(B2�01 f`2� O{RD|�scii��oload3�41%�ylJ�i�Guar�d$P�mP��k7�b]naPat�& 0N"�Cyc��0or�i���`iC00Data�@qug�c�3p[,`�3FRLOA�am�5<�3HMI� De�2(�1oc6�44�0PC�sePasswo�aA)qp��1p���{-+Pve�njCT���YELLOW BO�I� t�"ArcV0v�is���%���We{ld� cial�$_    �et�sOpA ;�41\\��5a 2��a��po0)@`@�aT1���5�0.2HT� @ xy��R:�82���`gp�P��xp�� 12�A�JPN ARCP�SU PR\A�T�Eh0OLwpSupg�fil5p�Q���^ l�cro�6 "AT�`�3ELdx�!���SSwpeetexn^$ J3�QSo��t� ssag�% 	T�eBP� ] !9M�Virt��39�V }h	`stdpn6����ro� SHAD~�pMOVE TF �MOS O � D�get_va�r fails ���ߐ  � D��E���� Hold �BustdCVIS� UPDATE �IR��CHMA �62�q�WELD}T�@S ) "��~�: R741-�kou
�b��m �BACKGROU�ND EDIT �Ò m41�0RE�PTCD CAN� CRASH F�RVRTO�Cra�.�s 2-D��r� �0r$FN�O NOT RE���RED � P�CVl�JO�P Q�UICK�OP �FLEN .pc��c���TIMQ�V3 ldm�PFP�LN: 燹 pl� 2���FMD D�EVICE AS�SERT WITg iC��sANġ�ACCESS M� �aŀo1Qu�i��<!�C"�US�BU@- t & rOemov��<�2� SMB NULAp�ܡ��FIXW��H�IN͑OL2�MO� OPTt�PPO�STwp��D��- �� �Add��adl. 	�io��$P:��Wu`.$ѠO��I�N��M��CP:f�ix CPMO-�046 issu5e�tJСO-|�2��130���SET� VARIABL�ESΐ�$O�3D �m�"view d�a`PWea�80b~. of FD ���u)��x OS-y1�p� h s v�D�5t��s ��lso �(� WAx���"3 CNT0 �T�S$Im�Z#c�a��PSPOT:�Wh�p��s�STY�܄At�pt�d?o GET_l���VMGR LO�0�REA�pC��M�`P�@ Y��0�EL�ECT��L��ING IMPR N����Rɰ̐sPRO�GRAM�RIP�E:STARTU�@AIN-��D��Q�ASCII�d�O�F L���!`PPT�TB: N��ML�Kdme�4��:�m�oW�all��R� �Nu�Qr� Angȅ��`d��thzo�n[� ch >`pܐ�r R2toun��H85@�iRCaylA�"Sign�0��pI,A�Thre�sh123�#.c��Hڰ : MS�G_P�єper �ࠡ��A�zerqo5P� A�  J�!fO�Imr � 2D�0�rc imm�`SgOME�s�ON�������0SREG:��^5� LB A�9�KANJIH�n�o��`c	��n 9dq�� -1o���INISITALIZATI��cwe��0= dr\ � f��aP���min�im90rec 1�lc0�:?!blem��ro��L�<3a �i� 09 ��b�d��w-� ݡ�0�w� uHQm@se�4SY�M��s���QЧ �090�Wlu� E�;BRe��jձ4�1����m ���Par��r@ G�Box f�o TME�ːR'WRI<���SY��k\k��F/�up��de-rela2Q�d��#5�betw�e�pIND��GigE snap��us5�spo Vn�TPD��DOs�~ġHANDL �`�Q�i�D��n�0 �f.v���Bop�erabil�` stmCQ��: H5@r�`l��L�
! ���m@ph�s U�IFL�PO>�FA�����ΑV7.��C[GT��pi�AsM��5pj�)@U��ine-RemarkO@�0 RM-�$ÔP�ATH SA̐L�OOS���v�`fi}g�GLA  �0d%���p��J� ki �q�ther�A� [Tr�`in�DW��4��2�7�� X�е�h��8`n;� C� R��:  6�d� y* it 35\k�wPay�a[2]_^�D1: g�s> �dowD2	SDIS�p�1�EMCHK �EXCE ֠�$M'F +  ��h�"��P��Վ�B0 c0e1Ȣ��me�� �c� !?��bP��� BUG��yB
:�@DŠPET��V0�0�T93X�XPAwNSI)�DIG��>��O  H5�P�CCRG ENC�CEMENT`�M�m�K 1A�H G?UNCHG OA�1�Tڐ����Sg\�d���10ORYL�EAK������L�C WRDN R���O�`j5`PO�S�PEްCG�V 7ont��VM�����W��@`GRI,@A�7��� �PMC gETH�0i�SUذ�>� H57�P0PENS!�N���ː� RE (i�RO�W<�³RMV ADD  II�=p���DC^ q�T3 A�LAӀ ��m��V�GN EARLY>���f n� ��衸E��ALAY7u�СPD�g�ˀH1SS8�OU#CH��D��Fh������PCDERROR�*PDE��� WRO���CURS�PٰI�p@N gҰ�?Q-�158Kwa���S�R �ġU3��\�aptp��@T�RF�@�R�\`�UB�U �`��#RB�0SY �RUNN���`10|�ఱBRKCT@q�ROq�Ԁ���CDA�X��Djj�EISS�Ucހ\��D��TS�I�aK�tXM�IP�SAFETY C�DECK "M6 ���dѤ�[`S U�)�8�4}P@QTWD��E��'QINV��D Z�O����a�sb_aBD�UAL@|�'QòFR��E�4l�6��P`?NDEX F�P�U,���SUF�rPk�Lb�ѳ�RRVO117 Ay�T��챤 ���FAL�BTP24�7���P?q�EHIG�PCC n��0�EoSNPX*PMM�QE ��)!SQ�"V���8T�bDC�BDETE�C��ds!Sˀ�BR�U/b63���s� 0C2"�t�s�'�!h� Z�T�7pS��"e���߆��,����߉ـ��0�
ա��ق�c�scr�ـ �dctrld.؁��$�fّ��!���qfـ*��878���-�% ��� rmґ�
�Q�R��78��RIـA�̑ (��~��Q.����ao�ـ\��a:P���a���I��ta 3 "K�:����<�#�o��t�p؁ "PLCF�"E!�ـ�plc�f���ـ-���maai�ـN���ovc���ـt�/�ـ����x��􁢐r674���Shape GeQnwـI��R,����ـT�іV� (5�ـ��II���� �`+��ـl���sga �4P� 4j�I�r)6ـŲ5=�5ѺI�n��ets6� " �PC���nga�GC�REѿ|�5��@�D�ATj���5ŝ�t.�!��5�a񯜳A�g�tpadb���Y�tput����������2ـ��5Ĺ���f��sl�q� 7�hexy��4����ώ2�keyy�ـ"�p1m������us9ߜ�gcـ����x+�H�a�j921��pl.Colly�����r�ВN��ڕr�3 ({�ـip����r��'���8�7=�7����tp�� "T�CLSj�|���cl�sk��D���s�kck���)�U����Ѱ�r�H���71a�-� KAREL U�se Sp�PFCTNj��7��a�a��� (��ѡ�� �ـ���ٹ�6�8=�8"�   �ـ 0�S�(V� �  lm� 6�9�9�~ F�)vmcwclmf�CLMl�0�`��60vet���cLM:����sp]�~�mc_mot����ـy���suX��60����joiT�J��_�logH��tr1c��ve%�� �����g�fin�der��Cent�er Fb!��M�5�20����g��  (�m)r,���fi ��1��a#z�� ��ـJ��$tq� "�FNDR����$e�tguid@�UID�ـ
?1��E7�q1nufl�60 �ـ>_z#ѯ 7A�x��(�2#���$fndr����c$���tcpS$]�CP �M� H�3ـ517��g�38�vC� gD�*Y=�F| Ց� ^ ����CtmgA4�P ��O�CG1ՑO7�Y��8�Etm �?�W�ـe�?�C�Rex��ے���Z��ڔXp�rm؁�_�D�_vars�_Z$M���V�h@����`�gG��ma|�w�Group�@�sk Excha�ng{@ـÖMAS�K H5�H5973 Ha�H5���`�6�`58�a9�a8��B�a4q2���b(�o#
k�/�غ`hp
8�0Y0/_цt�qTASKY_�r��pz�	h�Z�m@���������SDisplay�Im��v{Gـʑ8�OJq(P%���@xa���a�� ـ�lqvl "DQ#VL�t���q������Ϧ�y�����1av�rdq֏4ᩅsi1m���0��st��o���d���������v��0Z樁���"v�Ea�sy Norma�l Util(i�n4�|+11 J5C53��a�c���(���0��)�M�<�O�<� /k986TA8��#|�4�� "NOR�
`��1�_���|�su�� .������7���a!g�~y! menuu���g#M�����R57�7� 90 ̒J989��49�L�A0�(�ity�E�A�,`�P�m&��mh8��"8 2��܄����C�8_Sշ�n "MHMN�r%.Ը%� ��ͯ�s����i�Ը-at�Х_������֌ֶ��tm�?мz�1�����Q�2�Ͽ�z�3<zos�odst��
��mn�O��ens%u�Lm���hRaL��߃��huser!p�a����c~����Ը5�ɯ�����op�er���XԸdetbo`Ý~ ��L�UA��������dspweb���+�X�r��u<1��101W��הּ�2N�A�e�3!0A#0����4N�;2e�5��|����"��CalxN�0�O��Z� �0�O�$�S%j{�u���� 0S��}���ump��\b�bk968�!68�!��b�eq969B�9�%��F0b��? "BBOX�ۍ>�sched����setu~Xk��� ffH)�0��eq)��0�col(�1bxc��8�li�Љ�aI����W!i�e@m�rof$T�P EB!TA&@ry�|M427�*l!(T\�Q!RecX"H
�q�z�?$it%�?#сk7971�!71�{�F��$parecjo���A��?'����X�rail�@nag�e��~@]��D2E� �[0 (?:H͒V|x@@1ipMa���3�p�!�4�"4�u��3pa�xrmr "XRaM$��3�rf����ß1�1ꫝ0�yturbsp'G#��^@� �015: ��625t/~A��\BH�'ZD iy!:k�E�6�"A���H� �7��P�.��E!pd "TS�PD�}�T�GtsglD��kY��O�CiC�sRct%���Hvr�vQ���K�P,��A  q#-a�21�Y@AAgVM �r-b0 ��fdE`TUP h�im (J5�45 l) �i`6�16 V2VC�AM .CLwIO Y10k �5W` (F�`MS�C ���bPs��STYL�Sua28y kr�`NRE I��`SCHgRp�DCSU tps�h ORSR� �ua04��EIOCW`\fx��`542 LEX="�`ESET��ia,y`0shi`7y`"R?MASK�b�7o�-`OCO[�x��a7p3Sv q`t7p02kv6U`xv39_v�x�LCHRvOPLG��w03;uMHCR�3MpC�`YaP`�p66�.fia54; #��MpDSW�`588��ip1�a37 8/8 (Dr0c�5r94���r7 qj5r�5�5r^v�p5�"9PRST VR�FRDMC�Sx�a��-`930 �>�`NBA  g1�`HLB 3 (�a{SM�� Con�`�SPVC Lia2�0�#-`TCP a�ram\TM�IL r�PAC�C�TPTX �p��`TELN 96��0�r9/uUECK��1r�`UFRM setL�aOR ���`IPLKeCSX�C�pj�qCVVF� l F7�HTTP strbZ0zcp�CGy�8�AI�GUI�p7 ��PG�S Tool�`H?863 dj��q�M�Oq3
vJ684c�\$���sق��s'�1ےs�a96� TFADȑ65�1�Cq53 � oo�b1�44r-�k��r9�VAT��JO775 �R�6u�AWSMے�`CT�OP �q�`olld��a80;!diy�sXYY�0 e���i`885 '��`LP�`u"�`� 7H�`�LCMKP��pTS�S J%�
�W�CPE \dis�`�FVRC m��N}L�U002 
�{en%�6 65JrZ'�7[�U0�po��Ƞ�K���t� I�4 �URI�5�&�U02�2 nse�{�3� APFI�`{�4b�2�`-���alOP���1C�33O�͐t�ptsD`U040&g�43�ٲ4�۰j� "sw%�1`b�	�4�C	�5 ��w�x�57�eU061t��S�6ұrob9�15g�i��68����$!!��7�w�7�Ё�|%���"rkey��	3w��4?ǽ���T����8'�089�U#09���P��9:����2 &�l �9&�l2��9B�VrU15�P�NM� slA �3#H�}���1q�0v4ӽ7��108 	�eDэphc ��s�1�q�4+�1����A�5J/�tx�1����1]p!u�Qѡ�t�1������`��3����6��1�!p �`�о�- W�8�147 ase� C�U`sB�1 �82��1�4�8� (Wai��599 ��aU166�W��1�W�4� j U�6$�#U�7�3U�8�3�ȱ��B��1{��2 �act���6 "M#CR@�ِ4�1�������967ǑU1S93�3��6��2Y�dsP��2A��21���as�F���<�28-���E�2 wF���Q55�(��� ��cر5)�w���q��p����qf��L��$������q4d��2g�8q��8�51�""]�}�q��"< b������B]� � f�; `�̑ � ?8 16 (ݰ �BA��AAҰ�]���g :�!��`8 bbfo=� t� �j�� 7 \�� ]�� �2 �k_kv��74 0&!����W0H5���57&�579 h� L82 %"�\�4 3��5���5��1��59s4 U219 7,�-�6�p��6i�\t�chH6ur% �4>S3� 90� h��&�\j670��q���r!tD��4��&�t�sMg�lc�S�FrE�H��#F�����hk$�� sC� � ��"F�L��dflr��� �� ���fu!l%Z�gvPva���� sA����"D��3|��!creex�� �!�%�!�%�,���6�j6�s�!prs.�!�%�!5�hA�x�P 5�fsgn���/�/�,at<D�AD����qs`R svs�ch`@Q!Servwo S�!uleoCnA5SVS�!44�0��F��1 (�0A/ched�0,1�EA၍�� �2Q��0@��^�r0�U)1BBc��+� %P5)Q1�V�-#�3�1css "ACS�WVY88"gA@�`8!�/�0��@e���#M��C�3�tor�chm�0�- T�QMa�1�1M%'�9� J5lA598 *א1�!7)P8<P(1�̢A�ء%R1Qte,�!)E A5E`AS�v�� mLC6AR]C_� 1�4qc� �V�Ht!tc��A耥Q�4��R �F1 7T!2�S�EPBPQf-!�RtmkQ!p@60X��/�PRC8S�Q#�S�) P�2a96xAn`X�D.<bH5�1�U�}E� T�Qf#` aQ!<���F!�T!!�a4�3FcRO�Ttm�R!av`58�_�WP��MA$q�E88��>rp�in_��(�o�@e`AcB�rr��)u�!�U�etd�ѧ�U�Qovet�o�#$,�S�mmonitr42�=�Q�cF�st,"M_va�P`47M��V�0�! 5�8q���ameQ!Ɂ�rol�A��43�$Q0  Sp��1�0�1$P25�AKR  ��� 0S��(V�Ɂ)xj818\nl`mD��zN���r�MPTP"��O��qmocol �]/
�Y1�4Xa�@䁘�2�0i�53(1��T/ouch�!sؠ�2%qD2J5 !IU�٠��= b�0n��A�� ]�vP���z�EOWJ�th��Kwc���{��etth8!TH�SRXâm�t�o? "PGIOsRd�'z�wk� "WK�1�aL&MH�PH5�4�5�Q5�o��m`A��q@7z@6���1�8�a�PMor��tsn�@T�A�o�c���P"�����m�uA��T��p���T?��|�m4�TM�!2�5 4�>����m9�w�f�h�S�3G�qor�3���"641���8���Q!A�,HE!pR�U <�m�Re�h-g? "SVGN_��(�copy "CO�TA��U(��r#j0 "FSG��_�eh�j�f�@wA�SWwj|RbY=sgatu����!�;B�tp�AT�PD7��9 a790s����sg8!���GAT&o<Rc9  �Ħ�1�@t2`%1�&��1�bpv �1��&�1��B �1�8 6�1�chr��1�|v�1�sm��1�v����gtdmen�ps1�(v0!1��mkpdt�r1��]A1��pd��1�$&��1��mvbkup�.1��6�A��mk3un��G�pr���Gmkl1�e�P�s1��ni��0&1�ldv9r���glg�t��1��&���#�auth�.p�&��1�����) sud�1�7@� 1�G�1��\1�g b2�p�w 1�x6O�Ł4� 1��Ђ   946�"1����1�t\p�aic\p4k9471�wc��1��ictas-�Mpa�cck0m	8�	gen!1�I wl��Q� �stfq��q�wb���������vri/�4�^���B1�D��Pflo�w�@��Ac0ow�3<R50?���Q�TR�  (A0e T�0)B�Ԗ�cud!�0w�1��z�ac�$0�46 a� =�f�+p�aRa���!1�355Ţ1�F�ѡ�)a%|��;:afcald�� �&�0����%�f�m:�"�#�4�`��'a`"�3U���$��B1�! trac�k���@aine/Rail TrP̎�{(69�/�@ (L !iEYB�ʔ_ VB!Bu��a YB38P�48'7�	�F2���4��/�C�B1�3bŢ3�/�IUal��1�NT����VA��zQ�in�p�?0HVaen0�?DXWApuA�8�YqBzQtstd�0 U�@1GW ��]�j�VD����E&��VH@���o�peners^CO�`�ADev/w'~6�F8��񭁶��bA��aes�#1�]�ג��d����m�d1�k)9�@7�6��#1���/b�epaop`aO�PN�Wj�`��Krc#el}?�Exg���Y8`5Dv��tscx?tб�a�s FuvrCop /�Dw�nDh ��bAr5��QB�g�d�k�j!�� Pump v$Aᛑ�/�1�a;��M��T�q�i����t4U�1� 0�S��O \mh/plug�gr7G�h���u|bZ#��io�h#C{p��v(�ALI�O1�1�@7��93�Q51�91�����]4�� ST�
R��t�J989��/RL�SE�g1�@Cd�(M�1�/O�'�Q�)�D��G1 zq�H1�55'?��zq�tcwmio��MIO��$�tc�q"CL�01�UQcP�|�iEo��u~0%�l9� zp��v�1o���bQ�tzt����dtz�5I$��V%�rh#Inste�Q�� Co~PIo�qvRP1�hd�B554 (l�oBv��,�Q�H��Tcipc��oo�ڱp5�A�(
@��������"7`����aڰd�QCD �W�	����8��ڱ�rGcnd�_׳1p�a�ײ������Sb��a��O�2kz<�rpcrt�ᱯ�pٱdEc��S d��\���u�E!߳vr2k�pE A�-�x�_B�\"� choO�l"u�C��Y 1খ630 @ᗷ�@�� �ӿ�q�X�ԑ�GTX�? ��>�1chp "��XOh:�3�&�"5x!E��\p3 ���P��j�d 11�$h��Plo���ұ�c!h��3��s1��a�01���#Ar�� �0� !oCB��spq[`Jm:�k�7�)�vr�������a!X%-J�FR�AJ�Watpqrn�ev'�����fQ��D5��`��KrboT , �$��PG�[z!�sm�ICSP\Q�QP5y��!QP���j�H51�z�93QP7y�6���������5��R�6QP���NPR�`(�P@aam S`u��b��ĉa4tppr�g�p�B�	�Z�qratk932(q v輏�sc "iC8��~�atpr�_��qqz�;F�LGds�blflt{�ёs�able Fau`��CPav�aQ��~`aDSB (Dt$�t�d�A����QPh"@�E1��`f$*��3[S�� A�"tdj  "`PaV�Ohf$�1sbj!��1�"\:1gc��.��f%�du�550^CA�djust Po'int�b��J/��-��0�4�a昐A��j��O�N0\sg�4x��w�1\ada��O"ADJ�M�j0��etsham�SH�AP0���XDjpo  �e��G�a��UGQPG'(.��1:�k@ab5�J��KAR`�iagn/osti��!�a��66 J�C��a=P�(QL�Q&T�o�fkrldeP@���	  ��SQ��)�3/ρ[ypp��DBG2t�!O �U�Rѯ#��V��F( �шS7��Q�i�p{�M�ipper Op��Pq�����78 (MH G w�1Rlbk_�fTcBQ���0&�d038<B8�t��E��c�9_9�t��Tc��k����8 $q�SdrnpVǁ� �Qd�Ő6Tea�=����r Mat.Handlv �an`W�� MPLGv�A_�p�q(�sє�f����g ��b��a���f�� ����>@$w���� Dw��EI d���uu��m���fhnd �"F��  ��)���#� ��p���>��(Pa�0To�@�$V�!!�3#p��a�>��{�Q�k925B��26�q�3�{�p���2	ş�y���gse>0GS�qďėPR���T���a���t�p����{�dmon0_�q�Ŗ�ans���vr��{�=�����ͪX�<y��wsl� � pen��D��Y�WA��823X�Q
� G�0!'�&P��8QqI�Q�GQ �\sl ��!q��v����������֐�_�`����"S�EDGiOٳaQ�tdg�@T�AF8�F�� �BN���ÑQm�7���ڱA��g;Ж�Q���8��q�S�ileg�y�e���ϟ�9�F'QQ�<LaQQj517So�3-[JV�?�'�#4BA�49GA�WL�aw {�no�Qfԫo�H17D�#a������0t�  �>��LANG j�A5��5�5� gad5��C5�,TC5�jp .5�ce���5�ib=�5��#5���pa5��C5�W�~��j539.f5��]QRu5� Env�
5�5S��K�3y ��J9$5�.� ��;��G5�2D2�5�JS��p(K}�n-Tim��"���"¡�3H􅓹���\k}l5�UTIL"������r "QMG���,q5�C5��1 �"5�ړ5�s5�\kcmn��+��r5����utM�_�lre3ad���ex����"��\��l$"��1a35�rt[! -5� tuva��`_��5� �`CV����\�p ���Bp9t�box��_qcyscs}kRBTv�veriOP�TNv��l��e`��K���hg/>�agp.v1$�"�1$ptlit/DPND�BPm$d>n#te\cym$8$xo"��#mnu3�/�/�/�.5�/�/m$���UPDT it�e��.3 swtox95]�-4oolBD5 wb95��-4FR-4Y�� /2grd�-4��-4�b-4��w-4B-4.3 ��-4�-4'�-4�.3�B0l� /2bx "`�5�Q5I.3tl�7`��AE�#/2r l\�6��@O�-4 :4CoElD5eMa-4+�C�5�K�-4W�Q5ml�-4Chang95}�95�qQ5rcmdE�b�OZ��`6�5,r�7�6��70�5&r_+]22=_O]!2� c_u_3U4<_N^�57�_�_1UCCF�M�Ey��_accdau59#�6cAEX`� /2|�Da��4|aO/Jm�a�5�-4@�4�a AOSJ	Q�e�o�o�Y��-4��ZDQ-4sQk��?�@rtet�q�-4\$�3�q�eunc�.-4��4�q�5su�b�5��5E�q�5cce�@oRf^opm4E�o�fv�7�o�eT �c �o�nt$
Pte;�q �@�f\��k��6;��-4Ѓ -4�K�D��zh!-4xmoQv�b�q�et����f�"�tgeobd�t.���ƥ�etu � ɐ��ɐ��tɐٓ�xߟ�z��va�r'��xy&��pclJ�cɐ��ɐ��eɐgripsu����uti�����infpo��ܯ�B��ɐ������\�����ɐ�Ʊ�8�p��n ��ɐ%�ɐZ�mT���0ɐԶ��\�ogġ��p��%�p�\�palp�����s����ɐݵ���Ŵ����p�p����p�kagd�%�7�lclayY�k�A�ɐ��Adɐ5�p�������B��|�|�������q�����rdmͿ��r#inT�-�?�sO�Q߈c�̿޼s���ߧ�t�v�ߧ�h���s�tn[`��tX01�ɐ)�Dɐ� �Tu!l4�q��g�26Ϥ��upd����vr����נ1}�3�נ�ᜣϵ�il3C�U�l4����T�5e�w�s �ߘ�֠�߻�wcmx�(��xfer�~��tlk2pp���conv�朗ccnvݑ��5�ag, y�lct���n�yp��nit0���d���(��  ��ɐ 0S�(gV�U9al �#pm�Wse��2� ���V�C��(�z�@��A�0�|�m��`��&$��޷'#ro��@T/f(&���p1�mI� �,��$�+���/ �)G�?�+�� �L�ɰm ∡P?b6D�4 rg�������� ���?�9�� O�7�� ����>�/�T� a�8/�C�����E��b,֡)?�*��nq?_9�l�-!H�� � �HA |�p��QU1 p! �O���P ��S i	�Q�R@t�`�  ?���ɐ8� ��M�.Oreg.�ԃnO�o99� �� ���$�FEAT_IND�EX  �S �_��P�5`�ILECOMP �>���ba�Pa�RUcSETUP2 ?be�lb�  N� �aUc_AP2B�CK 1@bi � �)�R�o�o # %�o�o�Pe`�o )oe�oU�oy� �>�b�	��-� �Q�c��������� L��p�����;�ʏ _����$���H�ݟ �~����7�I�؟m� ���� ���ǯV��z� �!���E�ԯi�{�
� ��.�ÿտd������ ��*�S��w�ϛϭ� <���`���ߖ�+ߺ� O�a��υ�ߩ�8߶� ��n���'�9���]� �߁��"��F����� |����5���B�k��� �������T���x� ��C��gy��,�P��qi�`P�o 2�`*.cVR�H� *K�q�w��2PC���� FR6:D���/�T@` @/R/�=/|,C`/�/�*.F5�/�	��/ <�/$?�+STM D2M?X.��E?�=� iPe�ndant Pa'nel�?�+Hz?�?�j7�?�??-O�*GIF7OaOl5MO
OO�O�*JPG�O�Ol5�O��O�O5_�
ARGNAME.DT?_��o0\S__� ��T�_@_	PANE3L1�_�_%o0�_o�?�?�_2orog `oo/o�o�Z3�o�o@g�o�o�oH�Z4�zgh%7�KUT�PEINS.XML�o_:\���q�Custom T?oolbar(���PASSWOR�D��FRS:�\k�*� %Pa�ssword Config����� ���+��O�ޏs��� ���8�͟ߟn���� '���ȟ]�쟁��z� ��F�ۯj������5� įY�k��������B� T��x�Ϝ��C�ҿ g����ϝ�,���P��� �φ�ߪ�?�����u� ߙ�(ߒ���^��߂� �)��M���q��� ��6���Z�l����%� ���[��������� D���h�����3�� W������@� �v�/A�e ���*�N�r �/�=/�6/s// �/&/�/�/\/�/�/? '?�/K?�/o?�/?�? 4?�?X?�?�?�?#O�? GOYO�?}OO�O�OBO �OfO�O�O�O1_�OU_ �ON_�__�_>_�_�_ t_	o�_-o?o�_co�_ �oo(o�oLo�opo�o �o;�o_q � $��Z�~�� �I��m��f���2� ǏV������!���E� W��{�
���.�@�՟ d������/���S�� w������<�ѯ�Ơ��$FILE_D�GBCK 1@���ʠ��� ( �)
�SUMMARY.�DG篓�MD:��[���Dia�g Summar�y\�i�
CONSLOGQ�4�F���߿�n�Consol�e log�h��G�MEMCHEC�Kտ��J�c��M�emory Da�tad�l�� {)}O�HADOWY��>�P���t�Sha�dow Chan�ges��£-�?�)	FTPҿ?����C�n���mme?nt TBDl�l��0<�)ETHERNETaߑ�"������n�Ethe�rnet ��fi�guration���s�V�DCSVR�F`�F�X�q�t�%�6� verif�y allt�£1�p�1�DIFF�i�O�a���u�%��diff���"��6�1������{� ������	9�CHGDE�W�i���u�!�&��9�2������� ������GDM_qu�8.9FY3���� ����GDUgy/u��6/�UPDA�TES.U ;/���FRS:\S/�-�o�Updates� List�/��P�SRBWLD.C	M�/��"�/�/���PS_ROBOWEL��g�\?n?���? ���?�?W?�?{?O�? 	OFO�?jO�?{O�O/O �OSO�O�O�O_�OB_ T_�Ox__�_+_�_�_ a_�_�_o,o�_Po�_ to�oo�o9o�o�ooo �o(�o!^�o� ��G�k �� �6��Z�l����� ��C����y����� D�ӏh�������-� Q���������@�ϟ 9�v����)���Я_� �����*���N�ݯr� �����7�̿[�ſ� ��&ϵ�7�\�뿀�� �϶�E���i���ߟ� 4���X���Qߎ�߲� A�����w���0�B� ��f��ߊ��+���O� ��s������>���O��t�������$FI�LE_ PR� �����������MDON�LY 1@���� 
 �5�Y� 0}�=f/��� �O�s�> �bt�'�K ���/�:/L/� p/��/�/5/�/Y/�/  ?�/$?�/H?�/U?~? ?�?1?�?�?g?�?�?  O2O�?VO�?zO�OO��O?O�OcO�O
_��VISBCK������*.VD_[_�@�FR:\F_�^��@Vision� VD file �_�O�_�_�Oo�O)o �_:o_o�_�oo�o�o Ho�olo�o�o7�o [m(� �D� �z��3�E��i� ����.�ÏR���� �����A�ЏR�w�� ��*���џ`������𨟺�O���MR_G�RP 1A���L4�C4  B�9�	 �񝯯�����*u����RHB ��2� ��� ��� ���ݥ������ ���ި%�ߤA�5����_�J�K���J�8��I��U��@SF�5UQ�ƁQM���q� �E��Ge�A�F:�:�S��:1�?
]ޝ�@������ž�� F@ �%�1ŝ�J��N�Jk�H9��Hu��F!��/IP�s��?@�u��ÿ9�<9���896C'�6<,6\b����BhBs�S�B���B$��A�M�A���ʝ�A�|�A�ݰ�BI-AaJ4A7��0��$���9�A�?�M� �r�ߖ߁ߺߥ�O����AG�q@5��߯����4� �X�C�h��y����������BH9�� ������8�?C����F�X�5�
���P�X�P�s�`�w�����B����M�O@�33������\��UUU!U<��	>u.�?!���k�����=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!�� ۾G2kVD��@ D�� CϬ@�UC���Ώ�' �������-�/� C/�#/1��/Y�/�/ �/�/�/�/�/0??T? ??x?c?�?�?�?�?�? �?�?OO>O)ObOMO ��N�P�^O�OZO�O�O _�O+__(_a_L_�_ p_�_�_�_�_�_o�_ 'ooKoXi�Xo~o�o �oi��o�o=o�o�o BT;xc�� �������>� )�b�M���q������� ��ˏ���7�/{/ %/7/��[/��/ܟ��  ��$��H�3�X�~� i�����Ư���կ� ���D�/�h�S���w� �����O㿩�
ϥ�.� �R�=�v�a�sϬϗ� �ϻ�������(�N� 9�r�]ߖ�]o������ �߷o�{�$�J�5�n� U��y��������� ���4��D�j�U��� y��������������� 0T�-��Q�� u������ϟ5G P;t_���� ���//:/%/^/ I/�/m//�/�/�/�/  ?ǿ!?�?Z?E?~? i?�?�?�?�?�?�?�?  OODO/OhOSO�OwO �O�O�O�O��
__._ @_�d_�O�_s_�_�_ �_�_�_o�_o<o'o `oKo�ooo�o�o�o�o �o�o&J5n Yk�k}��� ��1��U���� y���ď���ӏ��� 0��@�f�Q���u��� ��ҟ������,�� P�?q�;?��[���ί ���ݯ��:�%�^� I�[��������ܿǿ  ���6��OZ�l�~� E_Oϴ��������� ��2��V�A�z�e�w� �ߛ��߿������� ,�R�=�v�a���� �������'�I�K� �7�9�?���o����� ������8#\G �k������ �"F1jUg �g������/� /B/-/f/Q/�/u/�/ �/�/�/�/?�/,?? P?;?t?�?MϪ?�?�? ���?Ok?(OOLO3O \O�OiO�O�O�O�O�O �O�O$__H_3_l_W_ �_{_�_�_�_�_�_o �_2oDo�eo/����o e��o���o��
%o. R=vas�� ������(�N� 9�r�]���������ޏ ɏ��׏8�ӏ\�G� ��k�������ڟş�� �"��F�1�C�|�g� ����į�?ԯ���� �?B���;�x�c����� ��ҿ�������>� )�b�M�_Ϙσϼϧ� ��������:�%�^� I߂�Io[o��o�ߣo �o��o3��oZ�u�~� i������������  ��D�/�h�S���w� ����������
��. ����'�s�� ����*N 9r]����� ��/ۯ8/J/\/n/ 5��/��/�/�/�/�/ ?�/ ?F?1?j?U?�? y?�?�?�?�?�?O�? 0OOTO?OxOcO�O�O��O�O���$FNO ����A��
F�0Q P T�1 �D|���@RM_�CHKTYP  ��@����@���@�QOMP_MsIN"P����NP��  X�@SS�B_CFG B��E ���{_��rS�_�_�ET�P_DEF_OW�  ��-R�XI�RCOM!P�_�$�GENOVRD_�DOCV���lT[HRCV deddo_ENB�_ `�RAVC_GRP� 1CdW�Q X �O�o�O�o�o�o�o�o &J1nUg �������"� 	�F�X�?�|�c����� ��֏������0�b�ROUp`I�HQP������R��8�?T쀟3�|��������  D�ڟl���@@�B�������o�4�g`S+MTmcJtm蕗�������AHOSTC�]R1KO�pP��a� M������0�  27�.0G�10�  e'�t���������b��ۿ����4�˿ų	�anonymous8�f�xϊϜϨ����л���%�'��[� 0�B�T�f�x�ǿ�߮� �����Ϗ�E��,�>� P�b������������ �����(�:���^� p��������������  $s����� �������K�  2DVh����� ����5GYk m7/�v/�/�/�/�/ �/�/??*?M/� �r?�?�?�?�	// -/OA?c/8OJO\OnO �O�/�O�O�O�O�OO M?_?4_F_X_j_�?_ �?�?�__%O�_oo 0oBo�Ofoxo�o�o�o �__!_�o,> �_�_�_��o��_� ���So(�:�L�^� p����o��ʏ܏�� �u�١ENT 1=LO� P!��E�  A�3�p�_� ��W���{�ܟ���ß �6���Z��~�A��� e�Ư�������� �� D��h�+�=���a�¿ ��濩�
�Ϳ�@�/� d�'ψ�KϬ�oϸϓ� �����*���N��r� 5ߖ�Y�k��ߏ��߳�����QUICCA0!����p�3�1q�M�_���3�2������!ROUTE�R�����`�!P�CJOGa�<�!�192.168�.0.10:��N�AME !"�!?ROBOT����S_CFG 1K�"� ��Auto-sta�rted`tFTPkH���s� �����$� '9\J���� ��Jv!3E/Y {1/b/t/�/�/g�/ �/�/�/?'/�/:?L? ^?p?�?�?Qcu�? ? OO/$O6OHOZO)? ~O�O�O�O�O�?kO�O _ _2_D_V_�?�?�? �_�O�_O�_�_
oo �O�_Rodovo�o�_�o ?o�o�o�og_y_ �_1�o��_��� ���o�&�8�J�m n��������ȏڏ) ;M_a�F��j�|� ��������֟���� /�ɟßT�f�x����� ����!�#��W�,� >�P�b�t�C������� ο�����(�:�L� ^ϭ���ѯ����� �� ��$�6��Z�l� ~ߐߢ���G��������� ���T_ERR� M��.�>�PDUSIZ   �^���U�>n�W�RD ?����  guest\��������������SCDMN�GRP 2N;X����p���\�KM� 	P01.14 8���   y���}�B    �;���� ����������������������~��\��������|��� � i  � � 
���ҕ������+��������
���l��.V؋�"��luop 
dy��������&�_GROU8�O.M� �	0�p��07�	QUPD � ��U��!T�Y�M�@�TT�P_AUTH 1�PM� <!i?Pendan�������!KAREL:*����KC�����VISION SCET� ://��� Q/?/i/��/{/�/�/��/�/�/"?�/>YC?TRL QM�P��v5��
��FF�F9E3.?��F�RS:DEFAU�LT�<FAN�UC Web S_erver�:
Y ���A<OO*O<ONO�`O<�WR_CON�FIG R<� ��?>�IDL_�CPU_PC�0��Bȩ��@�BH��EMIN�L���DGNR_IOG�|���S�@NPT_SI�M_DOV[T�PMODNTOL�V 3]_PRTY�)X�B�DOLNK 1SM����_�_�_��_�_�_o|RMAS�TEP&|R_O_gCFG"o4iUOD|Eo6bCYCLEdo�4d�0_ASG 19T<���
 o�o �o�o�o!3EW�i{���k�bN�UM{�Q��08`I�PCH�o58`RTRY_CN�0
RQ�6bSCRN>{�Q��U� 6ba`?bU�M��p����$J2�3_DSP_EN� M�ᆀOBP�ROC��LUMiJO�G�1V�@Q�8�?��{}?ŃPOSRE��~VKANJI_` d�
_H��V�W�L}6�h�1�C�CL_L��@�r�H�EYLO�GGINB`����Q�PLANGUA�GE �6�B��4 �>�LGW�X�f?�ҧ���x% �Ԛ�?��@���'0���`$�>MC�:\RSCH\0�0\�?�N_DISP YM�Ĩ�8|�z�<�LOCGR�B�Dz�DA�OGB?OOK Z�kR�`P�T�X���B�T�f�x�����������v6	�<�������_BUF/F 1[�]� I�2��H�S�h�d�n��� �Ͽ϶���������+� "�4�a�X�j�|ߎ߻������ߔ�ˀDCS� ]� =��;���C��5Y�k�}�|���IO 1^�kG t��� ��� ������� �2�D�X� h�z������������� ��
0@Rdxz��EPTM  GdR2���� 0BTfx��� ����//,/>/�)Ĩ SEV:���.�TYP���/0�/�/ �-�RS�0��|*�2�FL 1_��@��9�9?K?]?o?0�?�?�?�/TPѐ���"ݭNGNA�M��p�tU�UPSF��GI���E�A�_LOAD��G �%��%��_M�OV[�aO�DMAXUALRM�w��x {@AdQ:�<��C��
y@C��`��Oj�lM�@̀Ҁa�k �ZX�	�!�p+e���OΤ,RX_C_U_�_ 7�|_�_�_�_�_�_o o;o&o_oqoTo�o�o �o�o�o�o�o�o7 I,mX�t�� ����!��E�0� i�L�^�����Ï��� ��܏��A�$�6�w� b�������џ������ ����O�:�s�^��� ����ͯ���ԯ�'� �K�6�o���d������ɿ�GD_LDXD�ISA�0���ME�MO_AP�0E {?a+
 �  ѹ%�7�I�[�m�ϑ����y@ISC 1ba+ �����'T,� ��
ߺ�C�.�g�Nߋ� ��߬߀�����	�� �?���N�"���� �����b������;� &�_�F��������x� ������7��F �|���Z ���3W>{ ��p���/���_MSTR �ca-%SCD 1d͠�m/��/|/ �/�/�/�/�/?�/3? ?W?B?{?f?�?�?�? �?�?�?�?OOAO,O >OwObO�O�O�O�O�O �O�O__=_(_a_L_ �_p_�_�_�_�_�_o �_'ooKo6o[o�olo �o�o�o�o�o�o�o G2kV�z� ������1���U�@�y�/MKCF/G e--��<"�LTARM_��f���� �v������METP�U�n���5)N�DSP_CMNT������#�&  g-.a�v���y���#�_POSCF/�:��PRPM.� �PS�TOL 1h��4=@��<#�
��t� ��������/�q� S�e�������ݯ��ѯ ����I�+�=��i��#�SING_CH�K  ǟ$MODAQӃi��a���~��DEV 	K*�	MC:�HS�IZE�--ȹ�T�ASK %K*%�$1234567�89 V�hŷ�TR�IG 1jK+ �lK%%�a���  `������M#8�YP#����5$��EM_I�NF 1kڇ� `)AT&FV0E0���a�)I�E0V1�&A3&B1&D�2&S0&C1S�0=P�)ATZaߵߜ�H����p���	��A�9���]�D���� G߸�k�}ߏ� �����6�m�Z�l�� ��K������������  ������hs�-�� ���}���� @Rv);M_ ���+/*/�N/ 	/r/�/k/�/[m�/ ���&?8?�\?�/ �?;?E/�?q?�?�?�? O�/4O�/�/??�O A?�O�O�?�O�?_�O�_B_)_f_��ONIwTORJ�G ?���   	EX�EC1p��R2�X3��X4�X5�Xy��V7*�X8�X9p��R0B d�Rd�Rd�Rd�R d�Rd�Rd�Rdb�dbc2h2'h2�3h2?h2Kh2Wh2�ch2oh2{h2�h3�h3'h3�R��R_�GRP_SV 1��>ї�(q�� �M>E`Ѿ<H����4S�����>c'��@�_�DR&Λ�PL_N�AME !���p�!Defa�ult Pers�onality �(from FD�) ��RR2-q �1m)deX)dsh��q7�X dv�  ��$�6�H�Z�l�~� ������Ə؏����@ �2�D�V�h�t�2� ������Ο�����(�:���<��d�v��� ������Я�����t*��R,r 1r�y�հ\��, ������f� @D��  z�?���f�?x������A'�6z��ܿ��;�	l��	� �xJ԰�����˰� �< ���� ��IpK��K ��K=�*�J���J���JV尻�"όɱT��:�L�Ip@j�@T;fb�f�n���%�4���=�N�����I��g��a������*��*  �´  ��`�>��������n�?z����n��g�Jm���� 
߀ғ�%��Ī�9��� ��`�  P�}pQ}p�}p|  ��r�/׈�+�	'�� � ��I�� �  ���J�:�È����=�����6Ç��	�ВI  �n @
�+�l�$�l���9�A�7�N<�p|�  '��_����@2��@��i�f£�@��C��}C�pC�@ C���C��C��o�
��A�q� " W @���%
0�B�p*�A��2��`�o�R�n�Dz ��q��߁�������2���( �� -�����������o� ���!��o�M� �?�ff� ��/A�� ��v�7�a�:�
>��  P��2�(o��e�����ڳ�ڴD�?��o�x�"Ip<
6b<�߈;܍�<��ê<� <�#&�KNA둳���nO�?fff?��?&�3�@�.���J<?�`�M����.ɂ� ����lƴa2// V/A/z/e/�/�/�/�/0�/�/8�F�p�/ 4?�/X?�y?�K?�?~��E�� E��?G+� F���? �?�?O'OOKO6OoO.�BL��B�_0� ��OUO[��OcO_o? 5_�?\_�O�_�_�_�_�U
�h��V�W>�r_on_/oo,oeo�GA��d;����CRo�oNoD����A��o�o%5yķD���8C|�spC!H5"Z�d����a�q�@I�~N'�3�A�A�AR1�AO�^?�$��?��;��±
�=ç>�����3�W
=�#����{e��n�@������{�����<��~(��B�u��=�B0�������	��H�F��G���G���H�U`E����C�+���I#��I��HD��F��E���RC�j=z�
�I��@H��!H�( E<YD09ڏ�׏ ���4��X�C�|�g� y�����֟������ 	�B�T�?�x�c����� �����ϯ���>� )�b�M���q������� �˿��(��L�7� Iς�mϦϑ��ϵ��� ���$��H�3�l�W� ��{ߴߟ߱������ ��2��V�A�z��w� ��������������R��q(�q���������e���v����a3�8�������a4Mgs8������IB+����a���{� &&	fT�x��J�eP�P��A�O�	\���*<��R^p�����  ����*// N/</r/�)�O� ��/�/�%�Q�/�/�/p??'?9?  N?�l/�?�?�?�?�?�2� F�$�Gb	���A��@a�`rqC��C@�oTO�dq�~|KF� Dz@��� F�P DC��eO�O�I�cO��O�O__1_�c?̯��@@8Z^4R� � �� �n
 8_�_�_�_�_ �_�_oo+o=oOoaopso�o�zuQ ������1��$MS�KCFMAP  �R5� �`6uQqQ�n�cON�REL  ���a� �bEXCFENBw
�c�e q�FNC'tJOG_OVLIMwdp�rd�bKEYw�su�bRUNc|�su�bSFSPD�TY�p)vu�cSI�GNtT1MO�Teq�b_CE_GRP 1sR5�c\:�I�2�m� ��Di���a�Ώ��Ï ���(�ߏ�^���� ��K���o�ܟ�� ɟ�H���l�~�e����Y�Ưد�����F�`T�COM_CFG 1t�m�V8�J�\�}
�_ARC_$r��2yUAP_C�PL��6tNOCH�ECK ?�k �׸տ��� ��/�A�S�e�wω���ϭϿ������kNO_WAIT_L�wl�e�NT �u�kzw[5�_ERR!�s2v�i�� ��ߠ߲߾��c����^��T_MOc�wj�, �Ok�3���_PARAMd�x�k�tV#���=?��� =@345678901������ ������+�U�g�C�0����y��������t���UM_RSPACE�olV>H��$ODRDSP���v2xOFFSE?T_CART��y�DIS�yPEN_FILE� jq^��+�v�OPTION�_IO�YPWO_RK y'�5s x�fRuQ��82��2	 �	2���[ RG_D?SBL  R5s�x\�zRIEN�TTOp!C��oP�a.A[ UT_S/IM_D��b�b�[ V_ LCT �z?�*+^�)�_�PEXE�,&RA�T8 jv2u�p0"� UOP {.�PS0���/�/�/�/�)�$�O�2 �m)deX�)dh��X d��?-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O�H2
?�O�O�O�O�O@__1_C_U_%�<�O _�_�_�_�_�_�_�_�o!o3oEo�O� �O�v 1r(���(���07�,� �lp�` @oD�  �a?��cb�a?m�a%�D�cx�a���l;�	l�b�	 �x7J�`�o�u���` �< ��	p� �r��H�(��H3k7H�SM5G�22G���Gp
�������Yk|��C%R�>��qȋs�a|����*  ��3�4�p�p��pT����B_�����j%��t�q� )�/��aD�������6  U���P� Q� �� �|Б�������	�'� � ͂�I� �  {��i�=��������a	���I  �n @)� �mC���m��[�r�N���  '� 賔~q�pC�C�@D�s�pC���ҟ 5��
��=x@#�"7~9�^�n�B�I�qA��Q��� 0�q��bz比�������ȯ����( ?�� -݂*�`΁6���Am� �0r�x��m�lp �?�ffU ܫN�`��!��n�8m྿:̺>�  P�aզ(m������� q�c��d#?��m�x�A�n�<
6b<�߈;܍�<��ê<� <�#&1j�m�A0��c����n�?fff?�0�?&����@�.��J<?�`��l�����dѩ�e �ϟgߋ��d��Q�<� u�`ߙ߄߽ߨ����� ���)� �M�8�q����
��j���f�E��� E�0�G+� F������� �F��1�j�U���y�[bB��A��|����t�z� ��3��T��{�������t��h�y�u�w�>���*�N9K���A��Z�_�Cq�m<c��?��//(D///T)���pٞ��a�`CHT/A
$�x !�!@Iܝ��'�3A�A�A�R1AO�^??�$�?������±
=ç>�����3�W
=�#�>��+e��� ������{�����<��.�(�B�u���=B0�������	3�\*H��F�G���G���H�U`E����C�+�Y-I�#�I��H�D�F��E��RC�j=�>�
I��@H��!H�( E?<YD0X/�? O�?/OOSO>OwObO �O�O�O�O�O�O�O_ _=_(_a_s_^_�_�_ �_�_�_�_o�_ o9o $o]oHo�olo�o�o�o �o�o�o�o#G2 kVh����� ���1�C�.�g�R� ��v�����ӏ��Џ	� �-��Q�<�u�`��� ����ϟ���ޟ���;�&�8�q�\�(��3��,�����]��������p!3ǭ8���ӯp!4M�gs����IB+��+��a���{�E�E���s�����(Ϳ���Pe�P��(�{�4��I�[�իR}Ϗ��ϳ���,����  ���˿ I�7�m�[ߑ��H�  ߿������������"�4�F�X�  m�ߵ��������~�2 F�$�'Gb��ϲ��,��!C���@�s������ F� D�z/�� F�P D����������,>P��?���@@W
J}����������
 W�� ��&8J\�n����*� ����˨�1��$�PARAM_ME�NU ?q���  �DEFPULS�E�	WAIT�TMOUT+R�CV/ SH�ELL_WRK.�$CUR_STY�L G,OPT�]�]/PTBr/l"C�B/R_DECSN  ��,�/�/�/
?? ?)?R?M?_?q?�?�?�?�?�?�USE_PROG %�q%�?#O�3CCR ���6G_HOSoT !�!;DxO0JT�BO�C[OmA��C�O/K_TIMqE"�B�  �?GDEBUG�@���3GINP_FL'MSK�O(YT��9_�*UPGAUP \���g[CH6_'XTY+PE����?�? �_oo#o5o^oYoko }o�o�o�o�o�o�o�o 61CU~y� ������	���-�V�Q�c�u���*UW�ORD ?	{]�	RS��	P�NSW�V$ڂJO��!��TE�@�VT�RACECTL �1|q�� }��� �����4��DT Q�}q�c�(�D �  � p�t�t�V�v�Et�t���v�t�P��v�� v�t�t�P�v�N�v�!t�"t�Q#t�'�v�%t�&t��'t�(t�)t��7�0�� 6�� (�:�L�^� '�y���������p�Ӣ p�[�p�âp��Pv�� �v�� v�t�t�	�t�
t�t�t��t�t�t��@v�t�t�s���������@͟ߟ�����*��+į֯H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������	��-�?� Q�c�u������� �������+�=�O� a�s�l���������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_����_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
���_@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������0 BTfx���� ���,>P bt������ �//(/:/L/^/h!��$PGTRACELEN  g!�  ���f �|&_UP �~����!̳ �!� |!_C�FG �%�#f!�!��$� �/�/�;�"DEFSPD� ��,1�� ��| IN� TRLW ��-f 8�%�G1PE_CONF�I� ��%���!�$<LID��#��-�4GRP� 1��7�!��g!A ���&f�ff!A+33D��� D]� C�O� A@6B1�f �d�$I&I�1�0� 	 ?�"�+@OG ´yC[ODKB|@ �A�OmOO�O�O�Of!�>�T?�
5��O4_F^0_ =��=#�
K_�_G_ �_�_�_�_�_c_�_&o��_6o\oGo  Dz�c�of 
qo�oao�o �o�o�o0T? xcu������IK
V7.10�beta1�$  A�E/��ӻ�A f ,�?�!G�C�>��r+���0T���+�oBQ�c�A\i�PT�D;�{�p�"�B�������Ə؏�T�O'O�2�8�� \�G���k�������ڟ ş���"��F�1�V� |�g�����į���ӯ ���	�B�-�f��ov� ��K����������� �>�)�b�M�rϘσ���ϧ������=�F@ ��'�۫%W� ��W߉ߛߑ6������ ���%��I�4�m� X��|�������� ���3��W�B�{��� x������������� S~�w�8� �����+ O:s^���� ��
�<�//R�d�v� l/~/�ߥ/������� �/�#?5? ?Y?D?}? h?�?�?�?�?�?�?�? O
OCO.OgORO�O�O �O�O�O�O�O	_�O-_ ?_jc_u_$_�_�_�_ �_�_�_�_oo;o&o _oJo�ono�o�o�� (/�ob/P/&Xj �/��/�/�/�/��o ��3�E�0�i�T��� x�����Տ��ҏ��� /��S�>�w�b����� ��џ�������+�V_ O�a����p�����ͯ ���ܯ�'��K�6� o�Z����o�o�o޿ *<nD�rk�}� �����φ����� �
�C�U�@�y�dߝ� ���߬��������� ?�*�c�N��r��� �������0���;��� _�q�\����������� ������7"[F ����ο���� (�0^�Wi�Ϧ� ��v�r��/� ///S/e/P/�/t/�/ �/�/�/�/�/�/+?? O?:?s?^?�?�?�?�? �?�?�O'O�?KO6O oO�OlO�O�O�O�O�O �O_�O_G_2_k_� ���_�_�
o oJCoUo����o L_�o�o�o�o�o ?*cu`��� ������;�&� _�J���n�����ˏݏ O��7�"�[�F� ���|�����ٟğ�� �!���W��_�_�_ �����_�_ o���6b��$PLID_K�NOW_M  ~bd�j��#�SV �3e]=�:e�� z�����7�¿�������j�vmC�M_GRP� 1�P��`d�Jbd@I�߶B�_�
�_�����t��@� �Ͼ�^����ϮϪ�
� ����F��d�(�Zߠ� ^����ߔ߶����*� �� �f�$�L��Z�|� ��������,�>�#�+MR'É.�Tg��� 㢞������� ������������Q+ %7������ ����M'!3 �������Y�{ST'�1 1�3e�3 �i�0:o A >/g�</N/`/r/ �/�/�/�/�/�/�/? C?&?8?y?\?n?�?�?��?�?�?	O'2(.�:/j��<=O.3 'O9OKO]O!#4vO�O�O�O!#5�O�O�O�O�!#6_&_8_J_!#7 c_u_�_�_!#8�_�_��_�_!#MAD  �wd3#x`$PARNUM  ++q�5o"SCHOj ]e
�gpa�i=��eUPDpo�e�t>"_CMP_$�R`�ؠ`';�)tER�_CHK7u��0;�Or4F{RS|�2��#�_MOQ`��u_��be_RES_G' �+-O���H� ;�l�_�������Ə�� �ݏ����w&@�|�5��uu@R�q�v� �s�@�������sPП ����sbP�.�3��s �PN�m�r��s `����<���rV 1�P��^�b@cX��p�_$@cW�(��(�_@@cV�4���rTHR_INR|��Taud<�MASmSI� Z]�MNH��{�MON_QUEUE �.�bvg�U�g�bdN.pUrqqN��`{ΰENDб��EXE����`�BE��ڿ˳OPT�IO׷�{ΰPROGRAM %���%Ͱ믖o̲TA�SK_IQd@�OCFG ����o��^��DATAe���@�2�N�`� r߄ߒ�<ߵ������߀���!�3�E�W�
�IWNFOe�"ݘ�� ����������� )�;�M�_�q������� ��������n�z䍑"� !���OpDIT ���s�WERFL��#�RGADJ �&b
A��0�?���P��IORITY�av��MPDSQPX��U���v�OG$ _TG� �K���ETOE��1��b (!A�FD�E�p��!�tcp��!�ud��?!i�cm��FXY_����b���)�� *J/\/` ���G/�/k%w/�/�/�/ �/�/?�/2??V?h?�O?�?s?�?�?*�P�ORT3�Rc����u�_CART�REP�bk@SK�STA���zSSA�V���b
	25?00H863(�Ϩ�5D1�b`@�����s�O�O�G	P/URGE�B�	�yWF�@DO��$�ev�W�T�a�:WRU�P_DELAY ��bTR_HO�T{��%o�_TR_NORMAL{�x}_�_�VSEMI�_��_oCaQSKIP�1��u�Cx 	bO\o\@Jo�o�o�o jh�u�o�g�o�o	 �o?-Ou��_ �������;� )�_�q���I������� ݏ��Ǐ%��I�[� m�3�}�����ǟٟ��ͥ�$RBTIF|R�RCVTM.v+D�	�DCR1c�8lй�Cc��2C3fC6���?���>'�V;�F�em��%�����  ������o]����R�eo���o �<
6b<���;܍�>u.��?!<�&ǯ���)�ŰHB� T�f�x���������ҿ ������>�)�b� Mφ�qσϼϟ����� 5��(�:�L�^�p߂� �ߦ߸���������� ��6�!�Z�E�~��s� ����	������ �2� D�V�h�z��������� ������
��.R dG������ �*<N`r �o�����/ �&/	//\/��/�/ �/�/�/�/�/�/?"? 4?F?X?C/|?g?�?�? �?�?�?�?�?O0Os/ TOfOxO�O�O�O�O�O �O�O__,_OP_;_ t___�_�_�_�_�_�_ oGO(o:oLo^opo�o �o�o�o�o�o�o�_�_ $H3lW�� ���o�� �2� D�V�h�z��������ΈB�GN_ATC� 1�O� �AT&FV0E�0΋ATDP�/6/9/2/9��ATAΎ,�AT%G1%�B960�+�++3�,.�Hc�,�B�IO_TYPE'  ����Џ�REFPOS1 �1��� x��������?�P� ���6�������V�߯�z���� �9�Ǜ2 1�����$���� �ƿD�ё3 1� ^�p�����:�%�^�ܿS4 1�����Q��Ϻ���q�S5 1��ϚϬ���d�O�|���S6 1�߀/�A�{�������S7 1�����������y��0�S8 1�G�Y�k��#��G����SMASK 1���  
����e�'XNO��;�A������͑MOTE  ���ʔ��_CFG ������̒PL_�RANG���q��POWER ���^ ��SM_DRYPRG %���%��dTART� �V�
UME_PROs� ʔ�_EXEC_EN�B  =���GS�PD� #��4T3DB>PRM_P�MT_m�TQ �����OBOT_NA_ME ����׉OB_ORD_�NUM ?V���H863�  �t �ˀ!\<� � # 	r*!@̀"D|<���PC�_TIMEOUT�6 x��S232�
1�� L�TEACH PENDAN_ ����e����Ma�intenanc?e Cons�r���*"�/�KCLS/C� :���/�? No U�see��/U?�v#N�PO218��z��t!CH_L� 3���7�	�1�;?MAVAIL�a#����t!PACE�1 2�ٜ ��?%dH�9�eF%��<��L8�? H �9�O�?�O�O_�O (_#WTOfOxO�O8_�O �O�_�_�__o i� �4mT_f_x_�_�_�_ �_�o�o�oo .�5;A2@NROdovo �o6�o�o����4��I�N{3]o� ��S������ޏ 0�Q�8�f�N{4z��� ����p����8�@��M�n�U���N{5�� ����͟ߟ���%�4��U��j���r���N{6 ��Ưد����� �B� Q�r�5χϨϏϽ�N{7ѿ�������=� _�nߏ�Rߤ��߬���N{8�� ��$�6��� Z�|ߋ��o���������N{G ���� ���$
�� C�e#p��������� ����:hL���2��+��^�!dt Y�k�� ������� 8oR~q�� ����//=/ 7Ikm�/���/ �/�/??+?=?3/]?pW/i/�/�= `�� @NP�5<�?�/�) A�5�?1OCOI? #J$OVO�O�O�O~O�O �O_�O�O�O_^_ _ 2_D_v_�_�_�_�_�_ o$o�_�_
o<o~o@o�N<
O�oN{_MO�DE  +��iS �+��ox?v:A_��?'y�z	���o�CWORK_{AD�m<�q�/R  +������p_INTVA�L�`@�zR_O�PTION1� �u��VAT_G�RP 2�+�]�(���L��ԏ揥�
�� .�@���d�v���O�o ���dX�ß����ϟ 1�C�U�g�)������� ��ӯ�{�	��-�� �c�u���I�����Ͽ ��ϛ��;�M�_� !σϕϧϹ�{����� ��%�7���[�m�� Aߏߵ����ߛ���� !�3�E�W���{��� ��s����������/� A�S�e�w�������� ������+��O as���?�� ��'9K[�����e�$SC?AN_TIM�a���\��R �(�30(�L8z�_�p�p	
WtZ��2#Nq!»#Y�:.(/1��#M"2{$!!d��(~!�!�r #]) �0��/�/�/�r�)�/�  P5�0�2  8�?U?g?>1D��j?�?�? �?�?�?�?�?O#O5OpGO?Nq�%ROЌO�O[N![q;��o�t�Nqp]M�t��Di�t|!c{  � lM" Nq�A!
%�1_C_U_ g_y_�_�_�_�_�_�_ �_	oo-o?oQocouo �o�o�o�gS�o�o�o '9K]o� �������� #�5�G�Y��o�o�K�� ����Џ����*� <�N�`�r����������̟ޟ����1�  0�B|�_g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ�p���)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑ��ϐ����� ����0�B�T�f�x� ���������������,�>�P�J�V�   �1�������������� ��1CUgy �������	 �y3"HZ l~��������C&5/</+&��r! 5/q-	�1234567}8R���L{0�@�/�/�/�/�/?3,?>?P?b? t?�?�?�?�?�?�?' OO(O:OLO^OpO�O �O�O�O�O�?�O __ $_6_H_Z_l_~_�_�_ �_�O�_�_�_o o2o DoVohozo�o�_�o�o �o�o�o
.@R dv�o����� ���*�<�N�`�� ��������̏ޏ��� �&�8�g�\�n����� ����ȟڟ����"�+&s�C�U�:�Z���������Cz  �Bp   ����2/$@��$SC�R_GRP 1��(�e@(�l��� @� Z! �U!m�	 #�-�=�6�n�p� l�S�y(J�w�e�����7�3%Dʰ֠�o��ป���M-10iA 890�%90� Ɓ ?M61C �#�-�I���#�
\�l� ,�O'|�Z!�S�;�o�}�	n�����������X �,���Y" N�a����ߖ�i�@�.!�`/��m�����"��B�Š�J�H�a�H�9A֠p�  @. ��Dl��?���D�HŠ����H�F@ F�`�������;� &�K�q�\�������<퀈����������B���YD}h� ������
 CҾ?4#��0/v/�%���
������3�V�j�@���/7 B�*'���P���EL_DEFAULT  CԿ����X!MIPOWERFL  P�p%W"�} WFDOe& �p%��ERVENT? 1���I�n#�=�L!DUM�_EIP��(�j�!AF_INExd ?�!FT�/�7>�/[?!K߀? ��J?�?!RP?C_MAIN�?�8q��?�?�3VIS�?�9��??O!TP&2@PU6O�)d.O�O�!
PMON_POROXY�O�&ezO��ORB�O�-f�O#_!RDM_SR�r�*g_o_!RL(d�_�$h^_�_!
�0�M�O�,i�_o!?RLSYNCo.i�8�_So!ROS�/zl�4Bo�on? �o2S�o�o�o�o5 �oY }D�hz �����1�C�
��g�.���R����'ICE_KL ?%�+� (%SVCPRG1������D��3$�)��4L�DQ��5t�y��6�����7ğɟ�=��/�9��脆_A� ��i������>� ���f��끎�	�� ��1��ޟY����� �.����W�ѿ�� �����!��ϯI�� ��q������G��� �o���������� 9�;�翹�˂�ҏ� ����á������� � 9�$�]�H���~�� ����������#��5� Y�D�}�h��������� ������
C.g R�v����� 	�-QcN� r������/�)//M/��_DEV� �)�M{C:U(��]g$OUTYB`!x&c(?REC 1���` �  `  	� ` ` ` @` �!�!U+�#��U/�.�$`!�"?`!�)A8�+
 �P�b6 s�'��  �  �'� �    f���"�#�!U� ` /` �` ���=y �y �y ������` B� D��?O�%��|0��<S7  ��H� �0�_��? O�U` �4)` ��?S��`!y ��0�` �k� NPO�OOc�ʀ;[0�0�1o�  �=0i�O U!� � �` ` �,` �xO��y ��!�Dn� M�O]_�OKc��O�@�F��O�
__._@_R_d_If_�6r _�H�i@T_0�2�x�C�@��_��!r` �\4�P�#�_�fy �y �*y �y �` To�o�oh$0k �  �� �1   �i@=�o ;@�2�0� ` K`$|o��dy �y �y Dqΰ�! a�oh[�l��0k`�bR  Ȣ� lP
5�2` �Z` �(�c�4��Da��!��ta��;� L  "Ɣ3FG�ݢ �>` �`��� &` ` w��F��b�D֔DXb� >X��� �aĀ<Đ?g���?�?�?��?��ď"F �;/  #f�4���'�]W�  =� �� ���
` Q� ,��U�y �y �H��` !U|�b�t��"x1 �  �T�B�x�f������� ү������,��P� >�t���h�����ο�� ޿��(�
�8�^�L� ��pϦϔ����Ͼ� � ��$��4�Z�H�~�`� rߴߢ��������� � 2��V�D�f�h�z�� ��������
���.�� R�@�b���j������� ������*<` N�r�����%oV 1��, P 8�g@-p��*�P@P� }�(a*TY�PE�/e"HELL_CFG���&� �q66�0-RS�p ���//?/*/c/ N/�/r/�/�/�/�/�/@?�/)?8;�p:>����` %K?y?�?F=�J1J1�p�>�1�p)��a22!�d�?�?��HK 1�� �a�?AO<ONO`O�O�O �O�O�O�O�O�O__�&_8_a_\_n_�_|OMM ���_FTOV_ENO��nwOW_RE�G_UI�__IMWAIT�Rq�6k�OUTf iT�IMe��ZoV�AC�1o#a_UNI�T�S�fwMON_�ALIAS ?e~�Y ( he �o�o0��o] o��>���� ��#�5�G�Y�k�� ������ŏ׏����� �1�܏B�g�y����� H���ӟ���	���-� ?�Q�c�u� ������� ϯᯌ���)�;�� _�q�������R�˿ݿ ��Ͼ�7�I�[�m� �*ϣϵ����τ��� �!�3�E���i�{ߍ� �߱�\��������� ��A�S�e�w��4�� ���������+�=� O���s���������f� ����'��K] o�,����� �#5GY} ����p��/ /1/�U/g/y/�/6/ �/�/�/�/�/�/?-? ??Q?c??�?�?�?�? �?z?�?OO)O�?:O _OqO�O�O@O�O�O�O �O_�O%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3o�_Woio{o�o �oJo�o�o�o�o�c��$SMON_D�EFPRO ����4q� *SYS�TEM* . �"vRECALL �?}4y ( ��}!xyzrat�e 61=>de�sktop-b2�5t4o0:14744 ��q�q����yrw1}���2�D�V��w7cop�y md:pro�gram_1.t�p virt:\temp\�&��� ɏۏ�{|���1�C� U���������ӟ f�x�������?�Q�d� ������,���ϯb�t� �����;�M�_��� �(���˿ݿp���� ��7�I�[����$� ������l�~�����3� E�W�j����� ߱��� ��h�zόߞ�/�A�S� ����
��.������ v�����=�O����� ���*����������  ��9K]p� &���n��� 5GY���"����j;�frs�:orderfi�l.datmpback�//A/�S/f2�b:*.*	//�'/�/�/�/6o6x�:\}/� @�/��/<?N?�/7�%a�/?��?�?�?i {��?0OBOTO�?y OO`O�O�OeO�?�O �O�O>_P_�OuO_�_ +_�_�_a_�O�_o�_ :oLo^o��_'o�o �o�oo_�oo�o6H Z�_�o#��� ko}o�o�2�D�V�i �o����ԏg�y ������@�R���	� �-���П�u��� ��<�N���/���/ ��̯ޯq/������8��J�\�j��$SNP�X_ASG 1�������� P 0 �'%R[1]�@1.1`���?�j�%��ֿ����ݿ� 0��:�f�Iϊ�m�� �ϣ����������� P�3�Z߆�iߪߍߟ� ���������:��/� p�S�z�������  ���
�6��Z�=�O� ��s�������������  *V9z]o �����
�� @#JvY�}� ���/�*/// `/C/j/�/y/�/�/�/ �/�/�/&?	?J?-??? �?c?�?�?�?�?�?�? O�?OFO)OjOMO_O �O�O�O�O�O�O�O�O 0__:_f_I_�_m__ �_�_�_�_�_o�_o Po3oZo�oio�o�o�o �o�o�o�o:/ pSz�����  ��
�6��Z�=�O� ��s���Ə���͏ߏ  ��*�V�9�z�]�o� �������ɟ
�����@�#�J�v�Y�r�PA�RAM ��}�� �	�z��P��j�OF�T_KB_CFG�  ����ѤPI�N_SIM  �Ʀ�)�;�ɠr��RVQSTP_DSB �Ƣw������SR ��� G& ������Φ�TOP_ON_E_RR  ���~�PTN ���AݲRING_PRM�� ��VDT_G�RP 1����  	ʧ��\�nπ� �Ϥ϶���������%� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� w�t������������� ��=:L^p ������  $6HZl~� ������/ / 2/D/V/h/�/�/�/�/ �/�/�/�/
??.?U? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFomojo|o�o�o �o�o�o�o�o30�ѣVPRG_CO7UNT����N^rENB)�YuM�s�㤐_UPD 1}��8  
G �����'�"�4�F� o�j�|�������ď֏ ������G�B�T�f� ��������ןҟ��� ��,�>�g�b�t��� ������ί����� ?�:�L�^��������� Ͽʿܿ���$�6� _�Z�l�~ϧϢϴ��������VuYSDEBSUGhp�p���d�y��SP_PASS�huB?.�LOG� ��u�sr�����  ��q~��
MC:\Z�<
�[�_MPC`��uH�����q��� �q~��SAV �cݱ�ԛ�����S�V�TEM_TI�ME 1��{ U(�p+�t�����T1SVGUNS��piu'�u���A�SK_OPTIO�Nhp�u�q�q��BCCFG ��{�I� B��5�`5�;zC�l�W�i��� ������������2 D/hS�w�� ���
�.R@=va����� ���/��B/-/ f/Q/�/�/�� �/ �/�/�/�/ ??D?2? T?V?h?�?�?�?�?�? �?
O�?O@O.OdORO �OvO�O�O�O�O�O_ �H�_,_J_\_n_�O �_�_�_�_�_�_�_o �_4o"oXoFo|ojo�o �o�o�o�o�o�o B0Rxf��� ������>�,� b�_z�������ΏL� ����(��L�^�p� >���������ܟʟ� � �6�$�Z�H�~�l� ������دƯ��� � �D�2�T�V�h����� ¿x�ڿ�
��.Ϭ� R�@�bψ�vϬϾ��� ��������<�*�L� N�`ߖ߄ߺߨ����� ����8�&�\�J�� n����������� "�ؿ:�L�j�|���� ����������0 ��TBxf��� ����>, bPr����� �/�//(/^/L/ �/8��/�/�/�/�/l/ ? ?"?H?6?l?~?�? ^?�?�?�?�?�?�?O O OVODOzOhO�O�O �O�O�O�O�O_
_@_ ._d_R_t_v_�_�_�_ �_�/�_o*o<oNo�_ ro`o�o�o�o�o�o�o �o8&\Jl n������� "��2�X�F�|�j��� ��ď��ԏ֏��� B��_Z�l�������,� ҟ������,��J���$TBCSG_�GRP 2����  ��J� 
 ?�  u���q�����ϯ���˯��)�;�N�U��~\�d, �j��?J�	 HC���8�>����9�CL  B�m������z��β\)>��Y  A���3B�;��Bl�=��,�ɐ�Z�,��  �D	�{�F�`�j�C s��όϦϰ̖���@J��+�>�Q��.� |ߙ�d�v�����������J�	V3.�00m�	m61c��	*,�$�I�L;�D�>���J�(���� r�D�s�  #����D����N�JCFG ʖ�f� i��������������7�E��E�k�V� ��z������������� ��1U@yd� ������ ?*cN`��� ���m����/"/ �U/@/e/�/v/�/�/ �/�/�/	??-?�/Q? <?u?`?�?�?J�6��? ��?�?�?*OONO<O rO`O�O�O�O�O�O�O �O__8_&_H_J_\_ �_�_�_�_�_�_�_�_ o4o"oXoFo|o�o�� �o�obo�o�o�o B0fTv��� ~�����>�P� b�t�.���������̏ Ώ����:�(�^�L� ��p�������ܟʟ � �$��4�6�H�~�l� ����Ư���د�� � �o8�J�\����z��� �����Կ
���.�@� R�d�"ψ�vϬϚϼ� ��������<�*�`� N߄�rߨߖ߸ߺ��� ���&��J�8�n�\� ~����������� �� �"�4�j�X���|� ����n���������0 TBxf��� ����,P >t���d�� ��/(//L/:/p/ ^/�/�/�/�/�/�/�/ ? ?6?$?Z?H?j?�? ~?�?�?�?�?�?�?O O OVO��nO�O�O<O �O�O�O�O�O_
_@_ ._d_v_�_�_X_�_�_ �_�_�_o*o<o�_o ro`o�o�o�o�o�o�o �o8&\J� n������� "��F�4�V�|�j��� ��ď������O�$� �O��f�T���x����� ���ҟ��,���� b�P���t�����ί� ������(�^�L� ��p�����ʿ��ڿ � �$��H�6�l�Z�|� ~ϐ��ϴ�������� 2� �B�h�Vߌ��8� ����rߠ�����.�� R�@�v�d������ ���������N�`� r���>����������� �� J8n\ ������� �4"XFhj| ������/0/ ��H/Z/l//�/�/�/ �/�/�/�/??>?P? b?t?2?�?�?�?�?�?��>  @
C �
FO
B�$TB�JOP_GRP �2��5�?  ?�
G6B�=C�DL��0�xJ�@��
D@ �<� ��@�
D �@@UB	 �C��� �Fb  C��VGUAUA>��͘�E�E�I>��@�A��33=�CLް@fff?�@?�ffB�@Q�E-_8Wz�N��O>�nR�\)�O�@�U���;��hCY�@��  @�@UAB�  A�$_�_�S�U?C�  D�A�LwP�RO�z_�Sb���
:���Bl�P��P�D�Q�_So~
AAə�A�hc�ZQDXg�F�=q��e
o�@�p��b��Q�;�AȾ�@ٙ�@L�CD�	x`�`�o�ojo|o>�B�\u�oh�Qt�s�a@33@QV@C��@�`ew<�o>��D�u*��@� p�qP<{�	�Nr�@@�PZv_p� ���&�:�$�2�`� ��l�&���ʏ���� !�����@�Z�D�R������DT�
Fґ�E	�V3.00�Com61c�D*����DA
�� E�o�E��E���E�F���F!�F�8��FT�F�qe\F�NaF����F�^lF����F�:
F��)F��3G��G��G��G,I&��CH`�C�dT�DU�?D���D��DE(!/�E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[
�F���F��M�;'`;Q���8��`F�O����
F��Q��K�2DE�STPARS  ��8O@3CHRe�A�BLE 1�DK$.�
CP�%� ~ �
P�P�P�	GAP�	P�
P�P���
AUP�P�P�|�'RDI��NA���� ¿Կ���`�Oh�z�@�ϖϨϺ��΀�Sf�LC *ʍߟ߱����� ������/�A�S�e� w���������)M e�iߘ�$���1�C� ���%�7�IȀ�
�NUM  �5UNA�@@ ���[���_CFG ������A@6@IM?EBF_TTk���8LCx�5VERY�6�zK5R 1�DKO
 8�
B@2� �0/�  �� ����� 2 DVhz���� �/�
/S/./@/V/Hd/v/u_��b@L�
6@MI_CHA�NA L �#DB'GLVPCL5A�� ETHERADW ?�550�M���/�/N?0F� RO�UT_ !DJ!��4�?q<SNMAS�K*8LC;1255�.�5��?�?2DOOLOFS_DIk���%9ORQCTRL �mK���hM8WO�O�O�O�O�O �O�O
__._@_�|O�N_`_�_a�PE_D�ETAI8-JPON_SVOFF#O��SP_MON ��J�2�YSTRTCHK �DN�g?�RVTCOM�PAT�X53�T�PFPROG %DJ�%	qaRAM_1x7o�\APLAYl���Z_INST_M��0 �l�W�dUS8_WoibLCK�l�kQUICKME� �#ibSCRE@p}-:tps�@ib�a[p`y�"qp_uy���Ti9SR_GR�P 1�DI ؕ�0��z�@��5�#�Y�G��2  ����S��o����܏ǅ ����)��M�;�q� _�������˟���ݟ���7�%�G�m�	1234567�h����b�XZu1��{�
 �}ipn�l/ՠgen.htm�����*�<��R�Panel� setup@�}�6o��������ȿڿ o�e��$�6�H�Z� l�㿐�ϴ������� ��߅ϗ�D�V�h�z� �ߞ��C�9�����
� �.�@��d��߈�� �������Y�k��*� <�N�`�r������� ��������8�� \n����-�n�UALRM�`G {?DK
  � 	L?pc� ������//�6/�SEV  ��h&�ECF�G ��]�&��A��!   Bȣd
 7/�c-5�/�/�/ ??%?7?I?[?m??h�7t!�r��[ �3(ȏ�?B'Imf?wk�P(%*/O`
OCO.O gORO�OvO�O�O�O�O��O	_�O-_�<�d ��=�?;_I_?pHI�ST 1��Y  �(�  ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,��o�_�_oo ��9 �_�]936�_lo ~o�o�o1b�o�o�o�o %�oI[m ��2����� !��E�W�i�{����� ��@�Տ�����/� ��S�e�w����������L��QL������ 1�C�F�g�y������� ��P����	��-�?� ί�u���������Ͽ ^����)�;�M�ܿ qσϕϧϹ���Z�l� ��%�7�I�[���� �ߣߵ�����ğ֟� !�3�E�W�i�lߍ�� ��������v���/� A�S�e�w�������� ��������+=O as����� ��'9K]o ������� ����5/G/Y/k/}/�/ ��/�/�/�/�/?�/ 1?C?U?g?y?�?�?,? �?�?�?�?	OO�??O QOcOuO�O�O(O�O�O �O�O__)_�OM___ q_�_�_�_6_�_�_�_ oo%o/"/[omoo �o�o�o�_�o�o�o !3�o�oi{�� ��R����/� A��e�w��������� N�`�����+�=�O� ޏs���������͟\�����'�9�K�6o���$UI_PAN�EDATA 1�������  	�}]������ȯگ��� )  �$�ᔒ�O�a�s��� �����Ϳ����� '��K�2�oρ�hϥ�������������� Ha$�7�<�N�`� r߄ߖ��Ϻ�-����� ��&�8�J��n�U� ��y���������� "�	�F�-�j�|�c�������������� +=��a�߅� ����F� 9 ]oV�z� ����/�5/G/ ����}/�/�/�/�/�/ */�/n?1?C?U?g? y?�?�/�?�?�?�?�? 	O�?-OOQOcOJO�O nO�O�O�O�OT/f/_ )_;_M___q_�O�_�_ ?�_�_�_oo%o�_ Io0omoofo�o�o�o �o�o�o�o!3W >{�O _�_��� ���pA��_e�w� ��������&����܏ � �=�O�6�s�Z��� ~���͟���؟�'� ��]�o��������� 
�ۯN����#�5�G� Y�k�ү��v�����׿ �п���1�C�*�g� Nϋϝτ���4�F��� 	��-�?�Qߤ�u߇� ���߽��������l� )��M�_�F��j�� �����������7�0�[�����}�l��� ����������)��$ ��Pbt��� �����( L3p�i������ /(�����$�UI_PANEL�INK 1����  ��  ��}12�34567890 Y/k/}/�/�/�/�$�� W/�/�/??+?=?�/ a?s?�?�?�?�?S9S �*�=��U    �?O(O:OLO^O�?\1 O�O�O�O�O�O�O�O _(_:_L_^_p__~_ �_�_�_�_�_�_�_$o 6oHoZolo~oo�o�o �o�o�o�o�o
2D Vhz$���0��
�E0,/A� M�/�p�S�������ʏ ܏�� ��$�6��Z� l�O����<�?����� T!���1�C�U�g� Z3��������ǯٯ� z��!�3�E�W�i��< ��������C��ÿտ ����Ϥs5�G�Y� k�}Ϗϡ�0������� ���߮�C�U�g�y� �ߝ�,���������	� �-��Q�c�u��� ��:���������)� ��M�_�q��������� (�����~���7I ,mb���� ���3ƞ���� ՟w�������� /��,/>/P/b/t/�/ /�/�/�/�/�/?? ������^?p?�?�?�? �??��?�? OO$O6O HO�?lO~O�O�O�O�O UO�O�O_ _2_D_�O h_z_�_�_�_�_�_c_ �_
oo.o@oRo�_vo �o�o�o�o�o_o�o *<N`��� �������� 8�J�-�n���c����� ȏڏI��m"��F� X�j�|��������/֟ �����0���T�f� x�������?/?A?�o ��,�>�P�b��o�� ������ο�o��� (�:�L�^�p����Ϧ� ��������}��$�6� H�Z�l��ϐߢߴ��� �����ߋ� �2�D�V� h�z�	��������� ��g�.���R�d�G� ��k������������� ��<N1r�� ���;��& 8J=�n���� ��i�/"/4/F/ X/ǯٯ믠/�/�/�/ �/�/?�/0?B?T?f? x?�??�?�?�?�?�? O�?,O>OPObOtO�O �O'O�O�O�O�O__ �O:_L_^_p_�_�_#_ �_�_�_�_ oo$o�_ HoZolo~o�o�o��o �og�o�o 2V hK�o���� ����o�/�/�u���$UI_POSTYPE  �%� 	e������QUICKMEN  ��d������RESTORE� 1ݏ%?  ���,�>�b�m]������� ��Οq����(�:� ݟ^�p�������Q��� ůׯI��$�6�H�Z� ��~�������ƿؿ{� ��� �2�D��Q�c� u�翰��������ϛ� �.�@�R�d�߈ߚ� �߾���{υ����s� %�N�`�r���9�� ���������&�8�J� \�n��{�������� ����"��FXj |��C�������SCREր?�ۍu1s]c'�u2G3GU4G5G6G7Gy8G��USER)d.@T(IksQ��4�5�6�7�8���NDO_�CFG ޖ� � &� ��PDA�TE ��None V���SEUFRAME�  ��&!R�TOL_ABRT81/��H#ENBR/C(?GRP 1���Cz  A��# �!��/�/�/�/�/ 6!
??A*ՀUr(A!~a+MSK  u%4}1a+N.!%[�~2�%��?��VISCAND_MAXs5�I�](�0FAI�L_IMGs0`����#}(�0IMRE/GNUMs7
�;BgSIZs3&����,CONTMOiUQ u4��PE���c�� �@�~�"FR:\�?� � MC{:\RC\LOG�F7B@� !�?�O��A�O_�z �MCV�O�CU�D1*VEX3[��`�qF�"ᖉ�`(ޣ�=��͍_�� Z�_�_�_�_�_�_�_ oo,o>oPoboto�o��;PO64_9C��B ��n6�eK L!IA�j�h�aV��l�f@�g�o� =�	�hSZV�n�����gWAI�o�4S?TAT �+�!@�O���z$����5J!2DWP  ?��P G)����a�;@'��2_JMPERR 1㖋�
  ��2345?678901|��� ����ď��ɏ��� �B�5�f�Y�k����<N0MLOW{~�@�0ζ@_TIYH�'��0MPHASE � %���3SoHIFTO21"x[
 <���?\�� ;�a���q���Я���� �ݯ��N�%�7��� [�m�������ɿ�ٿ �8��!�n�E�����*	VSFT�1�cV�0M�� S�5�q� � ��E�A�  B8������� p�����ª��B ��ME$�u4�q���a{~&%���M��x[�p�30��$xpTDINEND]H^8t�Or0U?�ׄ[J��S�ߏ���s5����Gy�	��,���������ߍ�RELE �s/q�XOjFt�?_ACTIV��~8<��
 A �;}�<���RD�`��C!YBOX ������v��p2���>�190.0m.��83����'254�����`�� �q��robot�ę� ?  pHa�upc���u���p��r���ZWABC�#�-,u�  �r�5X?Q cu�����/@�0//)/f/�Z;D�q���